
module intosc (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
