// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:51:17 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UHCAONQQ4ojz0qiyEA+5xq4Fly9FMqcg+rxr3rpuB3YcLAWFeIRD4U4YUYYV+vm0
aArRgybPcXEVcdri8xliVj0dfW4vngrJlpTCduTagoVQSBweHLZMQe0J2KZUuf3N
uVuo2W4h/ZUpVgyA1tmz+H8/CWELd+322YSmK10ryt0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33584)
VEmKUmBGtOxXXIeOj4dHQL68/ReKqyjCEcs3v86Esu9LSLYnBijAbdPH92ed3HMn
mpfd6TbDJdwh/tNfyyhPyo6NWnY+FcaO53ZUq9cOpK10Dzmn94INGpFMHezRxCVl
9vSaL6wCk6LGMi8rsjjH/JWoP8XMEOKzoh9S3XFyFkaBXwHq0KBahabEiYDDbKm7
NzWXvAs1ei7j1XB27+4SSTIOYvvTE1+o+7+MlZ7kvrNSgydXNhVQntJrnM2f7TV/
/2B6gkMDqAytsxjXu57LbJw26J4HDPdJlVxSMZvOKGJEJxr68D7H9WbfTftHVgY1
2I71GPhoNMLneZaKUBmZTAoaahQfrSpo8o7hI/z6pXX/CMFLeytGhk9pCHrcRmdJ
ScT2XnB5IJRGixSGN0XXdf84V9GqmruQIckgzUq1Hw/82T6KyRBhVMr+vQgVUB0Q
F5d4BT9VU9rtqInJhfLBmxo7Kk/PUCgIRHXIfNB/lNJ/zWDFKxlFkW65Y9RIbwBH
uXRO1WEkAHe8UMcmVAAf6kBpWoKw027UwEReub01JgI6wqjUgn6PVDwqYzKBcONu
rGs6RPZR8ExkqyJcKHEC48BJ2f+lpAzLp81cxpvkTowm4zvjj/HsNtuBInuCVx7j
t07BiHYQ8sp15Lzftwls81ecKT58jhK89kgnYym4Wq1Q3adXkkZUXNX+on01oBPD
gahmcwNl5Hz8r47LIEqYyJGfJ4SZGlK31l9NvjX4vXxlV0lZq7+AyQ7QUj/i0gQe
1uDZuVCjxPX/PMuFs822gctOPnZjZPLbhB6+R01b3eI1mKTqaQLVBxvWa9ZfKe4/
KIKhM9fPURNFg5ZNnr3rVcrkT/pUUIAHapZTE9MEF2tsTgEqEpKazD+Vyy//6gYV
mKnrT9FjYl5K4jHn8SagZa5P1UeT7UvqlF2KUd0aVndhUkcCwmmkA00qLWeH71IE
bCs5jPyq3xSfIteKAIcTAJuthKjlcIdD4CZX1YkgoTXEmfai/odINcBDtu9T/Gcp
0hWjkMQSPvJvjlC8BXav/aDzI+NKR5uORxk69OX7EHd/iuyJhBf8tKVWZckRWrqO
/YlkL+JfTB2SOjV0YsTA5Acgd901ExBjUpBrWvhTCtWa3LZxBetikmyYFleLS/5O
AUxXDxhoqm1YQD4ogB+kS5XLnixMuSvbOHcWM5JpgirackOTEwDqStN6EjLW5C1k
qbX7NeOmksqHyVqvFBzUORCSMmFge22OJJIHzmDPAAK5yeWEVyA0d41UwPWQ3eqF
OTIzliTMK7ebEIra+UwAacrMBBOi+5KAM9vxRLOC4xTxtfC3cQ0ATwx7oysL17z7
gQNVU2RM8/o2KZNPi0hlyR3wRogZgybAMZK0sFhZ9AyhewDA6vJmOIAa2cA9BBcw
BJD3kfO6qfWMlD6orF4XKAaSDncwqUW02oumZAHW15M2ojDSr5zP4kM8XbIt15YC
8EzFRWC/XT04UroJwq8XJPIRryXqneZJkMp7l7lmf3m8NvrdabAILz9JWjbDwQno
F6nhuH+aQRBRemzip10UK9kaYDVuqoZ/vcXGQvEfeBpCc/8WA0w5Cf1sG86bA1FF
RH1Do6G3YyJaGmW9Jz7tCRZNmhPCiEeuPvVx1yPnu0k7ChTrxreZ4yyvVZc0uLGk
nAKS3AS+3t5nbOjSVM8/T922MuzaO0POSB6YYJcq+CI4fedNyHBFxvQPIjPH9Gn9
jZ1L0J8TH0RQzE7jutrP7Me1jvTXMdrCGmlC/dSF4mgDfX4wpIWFUoTpvdWrsmk6
U3t4gx3paGSr3bt+ZoKkM5Q74qkYz+JCxxvAlaJo1GdTdI/Oz7VkzSbs55iT01Kt
y4PGTOlSBO6f9v/HOOpx9RH+32TmYcLqLyYyzIbN8rnZTvLfOefDm0BMU/FEJn70
ZVFELhq7odk0sAVA257J/bbXF8VWf3Ub/kQzB746sLo5XDaM1A+tVuM7mNhZe7if
VEng0uDGaztuxtXE//IV/eEf3oPwf7UkWluKV3vnkY2xfC2ZZbAgik0k/Qbkf62Y
niCtzdlesE/mmGMlFgQZw7JMfEKBIUR+mo55cEDqQOgWUWZclnYhd5fX28KVwgnj
ypRgE59XA2tePmjV65B1QNrg15YX7I4VKM8zUKoFS9xB3Na0eJJ9kB/BXhOZ/52N
xEMnHhTrdCKavbJj+DGVdTPrHDDS+8eUcmH2jd7QXuHaMIsENeTyg0hwLZmlfUBp
qhf7xWh54FyizDiYWV8c5uJht45ckScfNYoMOhthmkmX8IGOgG15I6J/NBSxMXLk
72O6UG/JyguRF5NfspcCMS5szl5MDm0xY8XlIKyCZrSL3/aKlXi7bmI7S9gYIay1
bKugDWTuEky13fi7N7trqsUK5FgLfgKmpeELuKRnfZ9soPkzzny4J+PXRdnr6QiE
SYRJN2c346IRN6Ybw0jXUfQeteinaFecMbcI0gjvncxvQGfIJOrIOE/RJT48xAEk
gJIII+mIBgt8FF53IVHJkyRrNZ8nmUJYpvUgRo/PpACYLiZXw1mbDqibiX0wYtza
vjBMUzSVOxT+MwAmbSluDRgxo4ykZhj6rxHmaWxva1rLryF1wNRYUa2o0pRJroMw
3Ukz8JpA0XcPKIPAytO5XzKm7IO261DrLUhc9+h3S0RnKiIcgCS8CboilcFd3SUO
KA+/Yd4FIiguG8gMkLszHRp7w2OFStGaarEyramAqCnlsKuSyrSD3sfEaDz0ID31
FVuwz5HpmnSc+AXi1o4NbmLyoKlol1LBTxzGFHcJxYyUwRN0Xg2hZofawakghEMG
qjZ4l6TeEK53o/CRrI1fc4Z1LguvzkTaQlxUkhzhlNkjzKJfi4wIlfRDuAFcol/W
KvKt79gpd/8DWLtzM23ktxYLNEaAUytU3M7DtyV8RQeR84eTVtItznXngxXxT4La
sVKgn1Ln+jLkKalHPTV01xgvUZX4IE7TqfXJI1Hka6OTGTFIZhgExWcl+SCPiqIb
qnXmkekaWBvY63MXQAaCaNSvUdd0skDPbnKxpdC7vVZ8Ww1YC3crmPypCRlz5YvC
yJj59N42clHe6RN3rfbfarm7T7gosbVbfUMBRENdGMEgCjqbssuiXxDBOSapLCmL
nOnMtLzlM0jou56MsF3Ji07QGrwBAbBPOFjTYcD+x285mx/wRd2SkSAhbMnH9oQ9
yCtY9EC4OJZKrDMXxEasJ5QTSiiJrmf6ZWMsTc4bZfWHDEf21cUKaK7I5ilqyhfH
XhVFE5T6vebSEy6i4a78r7aLr2uVg302+AxG7EYfl/zI5Xf+0TWJ2v2wOX/TmMGo
BaQS468f+aTv0+7PRSJSsOflVxk3AgsWk49jy5Su6dlI4iTIspH53yVDxbFekmtT
KrY9S/K0sd9+CSm48Q05jmmS6TSwMdv7a+J/d9ExglroD6crcYD7iK30yeC3QPSb
inQuiYawDx3lffx6Yrxja2j/Ax2N1XI9CDgqc4wYGmEBh6s1ujJIaIORqA8FWpGM
vjlcEwR0dHNWzvOMu9G3LUs2foy7zl040TU8ZiDXVAJC7uqf4kZViYM3dp0SkxSx
05qij7CNSQjMNIttBpNSQqVrT03MPCa0bVb01AoBe/KjP0OKK2uvvhV0P+ZcLkHW
IP0XDlcUVvQfUCxGeoxHgww+45w0hGjiMLMZYKPadnXLRJ/G5ORrkWLPS+OGgHkG
3K7S/M+bxUOXZlPkUei/e80pww+n6hQeuCSq6KiGcx4+VX32lXaT0cwnTDPg96WM
hYN1xZ095zItnPndPh5I20voipWmk6MpGxTP6Vem3CRfEa1maUnQtskpRWXZJmTI
XjmozZV5kjobfreAOGeanejIDZioAJenjBScbY7Dv6I+8J/mA4scYe/MR2z6D+ui
RSBtqNNekhlMS/19A8ez9J/6PM19nTLeGq53lgbQxRW15D5v+Pgq78gcuC8jRmWr
tbZtNz4GsJDtZNrFE2Sd4h+ttKLeAWkotZnZKVLjHZqjpoLd8O6oyZ69rgDWX/5u
aEfolD/jEMymgdRd/V9MTKFLRa9dxyUBVxnwqKQigSpeln1dKfzUovejG+Se3i8J
lIIkzuHCQRjVW3uIN+o2l6s/oiFs8GMZyoSwtNI8+sFEFdo5T/4DhCkqRuEUnjz0
owHPNwW5Sd9TSThNN4/UGNz3L5+UICdw3/Rh6V2VJAe6RD5yIhpzyFWQUIrg45Hs
uBYgDD3DZ7H3WfwNUHKyWpeqaDb6hFO4IA/9PnmGvB5lfPA2WnMN/UUUMQRu7ogQ
p5HKRuoNHX4RJFj9S7q96148ofT4ONZCHcQgxt1eh8p63HNs3xeme63iFlzZddoC
lURBDplQsi0xGE4f+K+YkQMLQo2bChLtTIg9P1oxYkrE9c5oQlngy6yngQ8tOoqz
BdvTn0xQdnTj/ejuX/yxV64R2v5kEYOo/sIbbNUtcQXEabnnJqjMjnXFitvjFc7A
4/oPEf+XDTexvb8jVPEJ1TSqwXtAnWQvsNRHdM31Rz8ZxO+gq/3iNNB7dSVt+17T
rz5O5EZeTW4j/JMwkLO04I118fd1HyaVXKn7ng5wtn688zmwJdNUcurstMLX35oN
2nNWMcaGBRdIqB5+vSDgB9qCDNs4yf2yjVMCTPjq9hWOhfBSb6P8twkRTWhYey/Q
areeYkGonAKJKgMCtTQo06cGLaaEvcyUOYhjgQgWPG/dt+TuExkKKG/x9VRuowsc
nuz8+gV+bwmTVFQQgG1Y/Or4MJ8wLmmHm6ig++wRkcTg3cKpWFjn+Zj+LWldZMea
s585FSron0Xyy+totJqJo+tG0BvEi3gHL59aADRmVYdVt8NJYbqhvXwuvGrhVZjn
XJPceVJLB7GpL5OFYSk8AJtwtM+cZmu/2UJgHB7HBU4nhh1/wWifReET5KTjS0M2
8Pagt9yOTQfVtLAXBO33aI/vJrSC+4pFuHyzB5cSqd+IzX8sLfum49KwfPMtVLOA
c7shsTC8YG9g3kYD0FZbMCuFXe4WxQz022kw0VI1hhLVKupHJYVqCrcearoVlsPK
zwWBy9Zyko6cP09dJD8mzZX6gEnFbpoPHOrtNu5f22xgThogKeliec1NmPbFsFBw
oYW8bWRqoJNSuq6Amm7s5zGgaQGzKDW7K0jkZx/l9cKWK7reHWs68oQUPgWgoV9J
1mXHgsgc7E/AtJwolfotKBbiPOeDVLK09w6PuIKcOBpCtCkio28a5VIlTxpyRDjE
UjOKy9A5MhKaMM/Ru7AHUrjqFyyF00i04pze2DlYwkukD7dYo+t414/vGmJ2JLlx
ab6Dmc2hLXMzWSpSziw2MaY08fnu9xiszT89b2QhwsyPj8/+VC19aTej972kJDNS
Gfe9YVuCa070ahmXGjUhO6dAmmxsS1TXKl/T0DHdaK75b3Bmg6Cq4GRtsZ8MuvkU
kL7CP8qhK+aperMqTXz0yEi2o5cDk/6EkNCBM6eE8kWoeIhN9XjjHj3QMn2zfcSn
cgskGfhpslh++zQYN6Pcoms5hk2+cAmMiUYFtqhn2bcMAu496szs8/GnnjSFvwhO
McLqN66fsh9sLXgP8fHDqesTTXNbXKGA9MN5rpVjFAKbDXJqX5VwDvNTP6wBzeFl
m66/mEmLZ8qH5qIZErDKr3et2UJTfEffdXMSYTvSBZ77y81QVMC9lp//rAwHoxj5
Z1zxgx8BoKS7NXw1Rs+pDCVRMZY9j9YRRPvVp/NibInZmhlScGINcilWHnaHRF3R
YZL7PaYq1sI1i4bEtb37z3TgypjbijJECluOA/bbRHcqA6WqNZjT/Po3uLB/eIyK
n0oeVAfvrC6jj7XB5bJUuWES+jN8Ucr94jmpFWpjPNzuFFhYfpYQFc8om6jHPvOF
BrQYXgaoVwaHOA2TIStxlZ4adBh3FH9pF7KCiksjOV4NfvAaApsoJfKegz3euk6L
W4tNEiNpdcsn5yOL0ABTSiYbeamB1eA+D/G1EPjgV/mKEtZEBBiFoCTTtil8w5In
fVCZZgfWsDSajNsuoyKTRc86rfuCqmbqODdWjELrku7r5Eh6yM5Kj98UvAmRb9yk
F0E46ilLRs+VyjkkO74HGaw7yeLWn+ng9g/9z+ShdWFWnLMj88NtnhX4D0N4VCVq
uAHepVNmsspf/5P8D3gm3MugqJMy7eVTjnxHWLl15sfmFCqIP00Jyt4Y4owzPNXY
gE/XA7Ppp9eRDYRhEJqraPRJqwbVgwnSoprl20KzAaKC6QcjNWUlv6DR9g32xdMH
+9gBrOvF7rX+1nyFt4fj8wsGYyF8+jtWGA1stz/xlpeHe45m7qyfmoIz3Ir+3B38
9G5mN+BbBFWV2atZq1AHayWEdD61dVcH4+lQAgvlNzXva2EOHi/N6pEgsXPW+A1I
eEiEI9MwvLSSl10rweDIS/qVqbRnAHDYD0gtG9dPDK7sZGJiC+MkDRn16wcr/4Y0
JBDqeyJyuC4W4mZ23Kzm8Bmhn6nzp0I2EZDIxLMfCIKXgzy658DHGWtZUesxUKq2
4QF4jKCT9uk7z8KC4I9DXYN+qz8kvl66GxMb7t/rJKNIv7LR4w4NgZpta+MHkFgN
LkdziC1Wa5irv56kirPaOPgPSqhRD7QZefuCA5fh8AYq/vrjbi0qc17MmBoBWY21
4+GPfR5FCZnwuP9EQaKc1iNgWUlEkWWobXnG4DxwquZYM4+9Yikhfx8mxFq3ODVb
yS005lgnITl70FobzlDyifsN81HPKEraVPvr0cyOEr/oP/9jula76lWSHS3JdcnI
/5Xf7mJRN/MvevJbe1RjcjsJdmFA18zQKwWg6q9Vj76p4ZPO6jWpo3y/5g51QfUC
RoY7ZjcwxxQqVW10/Rh1yR6Yd72b9xeymLg8a0o8bSgknPAVxqB2IKn9JAFKcf+I
dnd1Sj2N8vFuebtY113N3A/9Btruha/oyqxu3NbbHzVC4klK3OHwv1xEmt/ZuWQ0
JQ4fe2uqwk1QkxoYt3cDLNZuPSp9VJmGsKkyuQzHvfJmQIDKpRGwIq5OXayUlphA
PnX9zrd2d5JnrFMYZcPrZyx0gtxuCRKcTpc9n0U7e6qumMRfgXoLe1QUFrHRDSnQ
nHA8XlE3658CEUIIS4payDx4/I9TlxxlSrLZAmeMz0Ot/PnHtec2x3cwVil5k9Qf
5+jVEbv2n/ALRkU2J3mzU9Dl3OIV+NAkwE/zH2A+K4sGeDFNfap6Y1r521geY9F+
P5jDe9vrfv4e0+G7xVAV6pT+ZociAmBUWh+VDLeMaqn1wWiqIcmsNkz6/TeZtL0x
cpyjILKTdJrnkSkwSdYti7v/oR7Wok6wVzs3eXpK/oJ1MmfE7qeSTPpiI5CmeHL7
VU6+qJ92CVv4SdqwZWfGMjHt1/Op9KXsBOR0x7gWy+tu6ZHd+8wwF/Eph/GPIyNv
QFBidzeTmtyY1CeHR2Amq/9PWwYOAgLNM/siFnRwjewihxB14qn2qAVFwXHZ85Gm
BEn/VQCaQ14Hl0MS+9E+Kw37/k0ZSDgTNGsss73KUwBjW5ILYv0Adso28EmnOvp8
s6aSVoXZ1qlNKpdtbJ6uN63e1qQxwN05Hary+m6OMTv+ORJjLwF3ZRCxFN6WV/0H
Kod5rm9licsb/cnYwkLLHZijsUtdR+FFy0gyKLdl5KjwVBVUIS3Dn9CpZ3y9DkE4
WROrxyPBhk7hDdXE8lQKQIFXrK97hPcDl+xX4lIMTTYDk45d3ioGX5p1UAdqV0fF
1pq99T8RPck+gBDEdsHjOBO0xbRkMZADob7h6My1U89QG1qDWg636s/9yt8Q46JV
2Z509yRoedzooY81bgLH52CoFLPf7inkQE/rxXz+EDDO9BWu+DBK6qrhozsx8hYF
Wk49ajYWJ+WBj46e5zeQCqQ1biB1FE2axafVMK07xaYTUPfuBCqmGLLg2U+L8bf9
EnaRDtnOSVJh9Duk9X9O3URv7wm2m8IRqW2AnTnN1CcNjCAV86ifeFyBHCcTRHlz
c00ELrrtWPbbf9W0OFm0gEd7PEWbrU8a0dd2Y8D/Y8pRlnbbtFRB+4IZ2NspHQA/
TdTQeFdeMuu+e/1NfC8TIH/zJ2ipSOblfp2QKH5t1ZPvkCaRIb5vTvm/ODOKy3dd
Pxyqll92gh+2WIBQyYAmWYLz2PYHMH0s5mkiC4c+dRl/rH1rx07K0aEQyRb4sMNF
jnJGv/Mn9zkGKDfy5UxauvpbajxM7ludJemx7C/H/gi1uIwHxrLp+2m8TxarJsqg
zi4yqgcUdDzrfbG/ysM+KICAE1ZMhnJGE4Ad/8Xml8+J/oT6oY110D6gYbvMatIp
D5/Ibg1AXWs0QMDDuDyPL/KiCUsI2aDE3u0b4NqTy8ncy1xh2CmvIuqvlFOJ8rmr
p0AnKvRg+qqVSQXYLsEbsi/xulebTCDaLAxodjkFBVvfFxVSnO62VaEoJZ8ITMFq
lLZW4qut3nXYiAkHrrHmsJygK6BqI5lyjviehS8aznr/ifqSRj1Wt12c5th2JTft
QB2IX9GI75shKWadDKyNggF+pAx305YT2QVmIRWmpNIwzdRtasiyQYsy9klqVUkf
mlN/ZppxCh8+1s2waZVPexSDbj9XdfZ5EtEauKmIHtrifLyegn9HBCcni8tV9lA6
wfSsQHAgMMVl0DTPsPX1PS+hCSdid6snKDqftz/KI7pQ8+COQvG3SjQoDqh0no84
Tfgd7jkgr/sPlLiXA5utbhhXQ0J/dCxWaBOor02qtnAFqAfiEuLPLVeaKZlDJYP7
49G+Uq0Tx46ZlTbckbReSGN+2+7G2Y+c/v31Qjh5CFQqjimBV68BKXM4ZGMW0LTN
OQyW2Uc4vQBbbidqrLvG7pL33AviWO9CL/F4DWa4turyvDiBZr4b66cslQVxXsFl
oJ3U4TX4hv2xY7oxCziVrN0DqXs0kxg35A+3Aaza7rPU8maoEiqvjLp1adKGqmSl
MsBq9VBdF0oweMxXVynz5FGYAIhVe3Plsy+aYUfUxZSA8VsSrtSDSiUlGtXO9KFr
ISdzk6oyq74JYjAxF3uVbJMqnoWJBe8QjQ7cVBqA3rGTgbt236pCZ7GtI+xjp8os
B14MiZZmsSNqnI6tSg7CaVNNGT0wMhBePcRrYukdAoSugmnu64SSMFPILdbv9WhW
qSzzaSgHpJKLSP6gF7Vae1+w1sziJTEU9+5cHP/V0s1bv93+Sj83gj4anOWE5jJw
NjyPPJh5CjGeFDeCobOG9NArFkj+RNxgyHwwavsbl1K5A83ieowM5iMTUFBVVj+o
RQlcxLKlDLzvvzolOBG7SWnuEBuHZ22ayzYlxbyu1XkXEYzy3n3x9hjbcezcuNf8
skUEeAjIVzPUDrzdEvzCANhctd72FKyA5s2tjhNnat62Qp/R3uuk0k/2g7RC+hio
mxdzz7c0aa66AqzhyQGQZNZ7WD+RxPu9KZIFaq8826YmEnOzsP/Y4a5q/B/azJA/
DKyvhpDbD6r0w0zb75rfy1NwKWBvdZKXoWlgICOmY8CMarvYGV3bz/WM688cPyYt
mgH31f8pm3sEs6uGmm5hQ7MGP7mZyO26gO89//hNAvbQncmkO6g11llfta/m1HGg
56iq85dxNOn0Oqs/0Ho9G9QB6DIRl0ICFkVVmRGdWcJEtRkRvoBJQX5FhiJ5tSam
MQ7EU828PJaknTvknWYL0OhKNAnvZ5SD94Z5jp5JnIxyX9eZsoPDQETd/LEUKajI
yRiZNlQp4r0KgrCsXSgCCpFiQOay4yUWZM6CR3uXaQ+NEZud8R/ztN2CQxodTlmU
ogl8yOsTEZo9TpNsKS2zFlcRHAF69B0WP9z/1dVRvUeSfofihgngJZClBtRzxZF0
Eq/oCdXaN+99on2L6SdeIgDaIG7ewWs7yCi/mOm3awvfint/bBqu+GfdLxq5QJob
0ukWTa04U+vzdFRpWSdCvUjLzOvRw2ZCXz0DueyjHVslowYtg8xIFwpNrBMxpr/n
0/PgX31+fTA/VJSC7z9C59cQ6hs9FbDP/mzaSzU7vATi5TMQPgAWcasFND0SXIWM
6uZwzMVv3XZWh3e1JXQLuPMaIoljioMnSqGgDp8TNK7BaydjkGp8lpuAEG+cn49T
5xt21NJ4EKS94dyy3xlppP4xK5+URUbotyZEnvepL6Zm9ZjfpYg6i/Mv/q57ZcrK
5Tk9Ket6ftQHXI+DKVPEslAFrxXH7hqOjQgQPI8jlXAYHLjUCD4aswSDLvxmYh9g
tbndIzkpO/MGJaf2bWTT9xQ2g1cw1rRSMQkFH6BQtMaM+muYovUjmtxHO2XROw52
y7EQQgNXyLJU1aAufniNqFt1Hr7Bqr/y9bExnSU2UEh+oICwBdSkwGJlsA0REdHj
P6KrFWdGMUpGQOJk9dAwFRTchTCkbI9VL+2sIS9CvSq1MbT9RCpADzk8S52uk5nb
ny6wcwUujdC+S9U69SnQMUTLRxB/zk8q5eEWqiRbDMYk74i15tOzQM14lSmaa81o
ijreMjf/XYH0DKA0OtNsiO5pEAoOvf7uJsKBUinBwgNX1wXtI6s5mq6ToDrKssE0
ahjpqxQK3JQwmuc+Owegd1J68VaZHZFDrpFfsmiCdPRvLOBHFg5FYgdX7weHV5S5
MXmQIewYfYmkXEkU6VWotHuC6e6CVmg8m9al8fBm+Ji2lvRJpfvYAOQwszFqSJ9k
kufRoipkc5ZvqN1NGHkjPTsN1R/al6yR8BBXJygfe1yW5IWPa/dFYSLZsAo6LvY9
biP/9pvvWQfeCBLHaQnHhxKtdJWroDcF8udhNzlLvY10yXN4FYfc1qpTPKGpYBO8
ArdKLf12N5ezX4uKrxUFRRxRKRSTu39ZmTOPjxMtge36xu99IInUOzipK84ot2F8
ozHd3nWXVjvu0cQSKG+alchE/vqPt7e0rBc91/SOXOKF4rBQDtI9u21mY+56JKU7
B8hrlAYMVVZ7pu/VtlvHeWFTi9lEIDqbJ9p04z4QmSYfXqHH6geznfO2Aoci0lxM
8oUxsH5wdO2Pc40R5wNEW6s45kP0jni5tS9HrHKYMwNHRwKNtTfN/TTgyoV84CUT
oCHBgHxis/sAVb3mczdFh+1TsTUu1336aNxNtCcMvXN1eRjyp8w87M/4V5U2v2ex
4fM9cMX7exbrUqDHQn1Ur9mvpV+qKC6hkHQVqHgBCiQdaVFPynlOsiGRb2pfx96H
AaRkaog2eG1rwh+bMfqVlbbLxcA0Uvadf3TaVkRwif0yTlF865sbk4fVuXF9Nq55
AhN11+hSuqKuwdHOnURkrXGZ2gnaLQZlbxh1YP/g1ZUlEuZOvaOZEMZ5T6YoeIBi
pdXkZ+jwGm0zpPydMz0OCgsOyVGb4T7qOM/I6s7XxM8OHv9l0OB8k8TgU01gzMsC
cLR1bN2pwBbD+icrh8G5khrywPW1z7rAJ0SKhRF3pHDytQOS9VVALU9lnCn66YE4
WL8qXSv0ZeMwYdqc3tVPLcNwT5XTaewm/0yDldtadcCeg/zqP+X/YrJrlLHA5caP
tkz4dWXQypeSZrgIWZvOL8enA+kxh6lo8TKGGqZYCRZTrzFrzKtf96/siB9Zp9OF
HeESt1qHyO0+z9EeaxxOuXYowVeEz7akAhm6IEL0/fKq+tTR2mj+n7whQZoGQp4g
okO9LMXzTmTlUIsBLmd3UWgOMCW1LOGG1nsQIpKRDbxNJps8jnCCK+/D8SNqVBKE
CefrWAznB+njNpd7Yf0VtwaoafxVis6S+qHgzibNOgJAY5bpnHw4CEeDza47yyXH
Xvf7G3LfGwvfcNOFKhhIX3sFUHCOyQAcfXiNKoh0QsDcr9HrF7AKQkDqlU79NlpW
AJXvx5LFnm/O5s2WisWc/lQHb0tGSJg7BGirIHWe6VmV3jqjRQh97iP/IOUOtiCF
453wT9n5v/FTzReBJIP/FomsHQ5JUsCNmtzJ/WX85vXbf+8ZUFiWUBbswybLoiLV
cui9lPvtJ+p5GEC1oUv6qI3qECue0XO70vfXwbQ0buKphFU4AhW/2eaHWxS9CQ+o
8YlSOklimabV6CorCa/gzKUIQAoJDjN4n5+unRc7+db8x2DcA8dL71XzwJDwMLUr
aJaSRSDhrG6qM1UsFoL+F1XzXHUE3LD+wSZBrZS8Xc2W3Dq1CP3hwVUHx2O1OQKT
cL+RuKvtjbeA6ISmUcfLKTVDdl7/E7mly7licXTz1tEK/7zT/prpPjWushffbT6R
rAz1UNE9qWY7fHLGN7/UBs66jJnH2Bk9/5fEz09KGltxvzzkr4++nF/X5CUpW6nD
/EsCWN9IONxB+VHUak7pneCsc5jE0Qf+2k/n8qUkIlJnVOmDtSkrC2R87PxcG9Z3
4SsBmpVX9wiQqJonyWkv/dy248iHTLMwGGUq9NvIHpbjTE4aKI7YJtaDieRG1Wuc
M9HX19hTGMyn72awM4KqY0H7u9Q0hmfLuagtjaDQy2MkjEyD24yvWxGAIj0PI2Ep
n4BG7tkiGUnDLMEb5f1Zy69KbRlBIfbnLuHQ8cMNlUbXTDJAGjgbiryEZTP+ujro
cKF84xFtGEcVwX7tH/iEtywraUPXNeHe/k12vYf1kfQxYg/vqp6uF5+Jw5nRVAt4
BaXBoVfnoNNhGWv4bHgNh8HaRHTRsJ0W7KkZ+W8xu3pfE/EIq6ifYoSIVclXsUtJ
jmnrvGNPBqCigBuLGvV92Hz0IIaxo2vFU3IN3t9zZiSqervKDMikKuXrhK2Irg3U
V6zRqC4KXwG+/dndyl+Z+PfpkDhvKm96N7+2P4VfkqFCwM/LpJ00Ia98fK/sw/8y
DMaj04JmYsCIgOxom/VsOy8+jLGTuDHMd7j6tdlf7Rkl/XgEJBiiXddQG9cEY0xj
8eZAtpITtbGg9UyL00WvHkUYoQhB7JcDA8m/ndXjVv2lAd5U4QpLT+8AXkHs80R8
B4yqkdchoFp0kcNIfwfNawrSRS5WOidUCLJxFc7YpHjhj7FxCbS1yUXP4Zt91qVT
AgTW87AXBSIRnqxXx6m3Ksk3FpKgd7O0tdsc1N8LAECnifYzPkBNHNgCVRbxcAmQ
JfFCFBEbJcQvR2aXq3lDDRY7bgXxYeeHkIa0MzDaLKsHccIpiAnsdOTwBELC33Nj
NHkeuRmlba5l35GPI5jgTmcLAmWjwm8tdBIgtewy9V3niPfiknR2Aoglq/Oz7PAN
an2DakXcRaWHY6kTcpx8d5m2PzZEhscmKbwz0NoJO5ow4T9y5BDVvLBGDJmhK/WI
q/TtuyJASG60NXOT8V/3hMSs0uAmYLewLBYWKsIlXTrjOHp2LNBF1wVBPHRLosEf
mbjPvMawrEVS7jSEXsqxI1xk63bRNZQNcMuxo9dxh9hnZ3Z1iiyTCfcGm145WS99
BvwllJzBNtGH52Hdm+z1vrkwB0O4dWznqPwGtd5bCKLNDNchmwJNCndWGuNiz8au
yj2MS90DIn1ip4iFs8PMKm+ooralWjHOIaCnLz+NzMuYdYpx+I+CqflEkBdAZw8Z
R7zGqloP2xFwskAUHU0eiTEVcKVSwjyeJn1Yfwfrya+SCouXKlmEDEuEnDu/YiJ4
6HZIWgdzlQ3jpFAONnUapXtH17B0U3g3hQwQ+CeWVz4Oy8yc5woXGipg5aBh+zoA
CrTSKGFexJ82nSwMRufa/cephI3wWetvPlNmJGxrOXt68SQ9glhMuF9SQenm9fr0
k8kE9gSjpIs3/S1US1duUhlHBSHUBFp8PWh0J41jmcSyspLGRFGypgpuYyxVo8YZ
e8YETaQHsLAyGmvy5SvnpHFTJ9PezVn0ugtg9vSOyy3mzJfAqRBozzeS7znk+K9S
eACOLuwnXDod3qRuynXerAzj4DQjBS+vgYq4Ryw67qwuvcsf4Cx53kcMAWJjuZyt
QFp8cjwI4ovr3/V9lNlFangdKzXUOQxyoWKr9xyTJt082kD9m7ACQ9yrpuyw3VlJ
zyfG22cdRncTCcBg3antWWusMd6KTaT235YZRwGfzpjV5ZsTYW0PJIoQNckvUgs6
5q4AHL3vhXAGeU+B3PFyw6mgs4wCu3P1AJZfXrfyObOGgXIvBK7L1r7EoyiJWFiY
csituJB7/vFFetNU6bHH9rRc7M7c011BA7HMzvTatU2nNIThebfyzGg+n3sc4QpT
6e7lsx7mBpiPs9QgVP72OGUklk5D2qiHGIi3tIlMuPKc0aIRQoIJbg1xhvqeY4Ew
hJvNE4o3lKuurP4JfWWTI/nuQABtoBy6FEfNl+tdhlb8Bi6KLnnwP+ZdUrD6tpH7
wh/+UqDbI2LAk51va4k6VU0geG85gBNA7cJ98jbWdJ51P/2si2ksd9GkO2xI58qD
zO/JtHr0GHe0EmImEJG1/XxkO1Qm/KhUusEw3/OY7nf1j3DciOVJedBg8J5QAE6q
JOl8/9zoP7Q7PTupRHfWiIslaaZsXdO1hM1Q/7N4kTaOhR+kuG7AM0khHuHmyf+O
Y0NLDjRswr5AoU62+4KYEHN+Y5G2PqbslckyzyeAOgL1F+PozjJncpgB89Vw/Bvn
bqH/imMVbZmrkuw7+GPaeH/uRSpvseqUolzHlpVxWAwx4XYsdfMWaiiIJKUVZn++
srKAKpmSgjkS4bKDHkOIp6la8zXSB1DgMFDbyszKimKjKRCzqzZgEq+grkeOrCAv
cY4Sx6SZsx1OUQ4fhJx1NCDQQ00Z1eB+VTsDf+sQoxHrVuTSOvruesYzOk04Arxx
MTwihUu2NImLkzRM6ASg08xXeEzUdIlYA7mS/c6YmNj0hClLRLPF9Ep/jrXnCr8N
aY2ZuUU/oQOS2f+cG3fiM0xAmrgLhhIigV3TCepZRyfn2hJeV6Plrh57n4sM0qE8
LpcZtqbygcW8rw0mXvAaB8EZ2C5FV4IqTeNnC9jDz+tFrUoUCe44zgM7pSGMJXFg
GVlYmsyTSxQ/cRCHRegOYA6HoWGfpOunR2Xlm6KMSbeVBI6NbMwES+A2eVspAlzw
8zlOzc298T0y4rVGG1kKBIkKLT4pXS9BvHodFD9gaAlhOFY0KrsTB/vv8Hj/oai2
2O5A/r90VGGAlEvuRIJ/jK73+YZ3TCPDBN5oODjTkKW0NA2tuHvPBk87Da9RxGR7
yGGpYuzabwnZUQkeECMf3FjKkRxNu2ChByNdmtEl9u0Q1xYXTBV7NQ1HI9xo/Qzd
+cvhI0m36W6mt4jW++EGa0d3WmtzygNeuANaaSe3nTgNOWYRRbGcLFFHj9mWC3Hs
F+Svfk7vrZTEV2zzcTtoyWifllk0nx/f6iHUrr6Q5D5RIViltBnjm4YRuHFpuO3q
b12pofi5hF7rg7T7OKMZL9EK1+BXyPWkqnzFfurJBC5p8v480R2avVFlSScJaukT
wL/IOO73HcpwHijNukp74uHj3gYpdg4A5uYRlUV4sN6rNoN2h4XBPWPbutUo3VI2
ym+wmWnqFaQcTWfa11ACNMCSCwJ57cXZAQGVWVwKTVuylOUcgpEzCnOj8CvFqKVF
moIOIBIoBiDaF1vxIjVaPSzMC5MQ2JuxohJ9o6OjsIMTe7qmClcobqd7eovHRUSH
F9CMxVsPDVCcc6mfdlbCQ/26QjlMTGqKvMPQhu6jKyamuRnQHUJGWkTxpvGg5kv7
Mpg6L0/lCuYQXHUIbUUn8Bk2SBsrZGRWAONtp1iqSZLOoMihO5xHwrCF17pwr9kr
WiqQTRC0/0ElCKAvnCesAkVmBVsKihRMaeQZBDdYWG27qMKQX8wtb4qHfSBh+Gtc
oynBRJZ/KLBDej4cGieDhrwB0qD3ONaqxcOAxjzw4oD8ZZwa11d84BtNoYeK1gTJ
6D3ObRAnkQl4P+EU2vVjtz3xYvFT7wwHDv7ON+YYs4B8T79jSkmcuLAJ46t+g94P
gPq6w82aoe4+SuOIKPgLGcQQm8yXOE2ffNdGoJsZ5Tn7qZLBX4k+iWbnmecfe+F/
FF8cqmh6ss2DGHmCDAv+yqtDQYY2KfFLcRxWG3ygtwCanw2tJb5+aMSrGi5bWRK/
roSi+DMwpZ/zYfw5UDI9zxhaqRMBtA3IQoqy3yaW2JianrxZYQeYpmqme1b/7+w3
PhdorEFpyXcMs+aRRXEhlqw8e2owOH/2B4apqCyGLWfHIgcHN8c9okCFRB/UHfDm
s75Px5kKOy9CMAwh4CW5ug25dN6iGCToIL8jRNFknvE+4qBbALTBUYxOjP3qyHDZ
4t6eYEQ5xSsKlTUgflRl5Kez69Hkc9kc1sC9S70dwXiGA/PE90dyhbZmytJxba1q
PJEstGBp42uuApr95FqGKWV3JDmy20oDWIhpoTvwG9Q0icW6bJjJEwIIW4rPwu0s
EtGCXiUcqVctTaKHjzTm/T8xP1L7Hn9NGHA+bb4ufCaCQHx6F0m1+HCEHXTh8vxr
GXtt9PTkFCvPy09c85qmGs4zNl7lYh04o0GwNfjd/IcND817Z7O7kX1IyHk8NpfH
4TaOJ5Zb6vvAYRY+W88Jyt1XpqF4XKq7OQA0PBIhFcKnMJRLVcGUgzplrRCZhRBN
vB6qbY/pD7AVmXQxRxYEVM63bo2GzhaheePzbsB8k30lsfXT1a2onaaja534M1Sd
Va9q8LxG7Dcw1XbdJc9ZRMCuAKbJXwMv8DDD9Q2lOJnGq2+9dofZbXYteGzO99w7
8iVfH5jru1j4tXp8ukyjAL0i09b+zTm2f/zop1UXR/j8MzrN8vG25fkVM40sKb+X
OJNVg5EHvwRYc4bu7rqIbSybhN1qlGT3u8/PhF07JCJ9j9NpJ001yUVBCczXjFCx
eFIh9gf5kolstKSQ5yTCHXb3+RL2cQSdBNfVbRF3LjOyTgnCTM6ajtId7zYZ2lZw
zXowg0otwk/urj7rODv9fgM/lNU/J+BZC8WbLv9Ji2RsKmN8+4ArmD1GZjsZRBnu
tELbHHRyYPfPQeZdbGdq/847/uKZtOOH8cnX92/lNxaR/cnjNTRX5/6qeNmM/I0p
iqu1gMVSSBFI9kAiNDUY0LTJLxll/CM3Qe4JpulVvJm2isM91wyjrwI2a+BnBA8+
pK0CNTC9obeKEiqW0xZdlufrvIvlQSC9NeFXyxBlMif1MpiWyHe6PbGaJUrmL2wx
40hdNjpz6hNdjl+N3SSkS4tpISQS7AguaMe6ig+6y3praSsqW6UwZDLsW2EiCY1w
fUdxSX3FVPFCaiYlJOZxuqCUV44WdEzvVT5kMJ+CF0SdPbleKNSVY/an5QThk9+x
QZDy9Cm9hlJWlbvFq1/Mvqq0moQ9gzibksPHaQE9JVP9CJkI8R3QYddb4nOWLbtI
SV/WKiWdnB2iMu477Wj/VLnXTP58aTBgJm63XRCT6mpA7dQ6GFSIEmT3ssqZEQh1
VEeQvX0tnO6sV0jJDkYvqH5zy4BK8RDqGTIh+E3/zr8ZyFOGnoCyQc5eUh4hONuP
+eOc/jEPG17yxaGt91hkb780lAiTMzegm9+ECwFqjcLKIhXf8PWdELL4GYWSUWX6
Nu7ozaMwntyEoYYR68WlTwjIxflaYaaZH1Oy0ncoSwDW9BAI7Ip+BbVhZeabHOaY
g3SH9efmWuaMpleMnB3w4lUbRnfL1JMCxcP/pzNVosn7Oc2imaS60HNTGfJ+a/WP
nlDXrzKYbdIKyt3Ooel27lkX+kL8gmEKnRHrNsJoKkntj5b/UL1CL2aIKvLfkxL8
pGbix38e42A9dI1PTbUvQhgmCI5VhxH9uJIDfyQ/UQz6FdPjH6ttOl/H9ep6iZBp
U0bIRssTUJ1yhMGY93liWhBStlML17CVoE4cWBQbVpgNgkOjOwWlojiBHKsHkouG
TnROqoSFoqHEN7syRoYxGUzi5Nbli53so0oz3cZq3sex3XfFjV0HofLu7v+icS24
gU8dOT2VUmKKy23UtZ2M+/fmCol6AWSZLm82Bn9Kme7ww5WN17nPVUT7WodOl4Du
OpGmJY1/pH91gwf1MvP66yzhYHJla6MAxpyOiv4OKmiauKBAV/GFn3BxWGsFhLft
XyzYk36zSF7c7l33YnslJhkZCDN4/I26DQ7pHXeYFPyhYlC7JozXC9mW4fHm5gp0
n5UKHjboSqya9b5KtyRN/d+05T46HVLKpN/rSTFes5G/MkgNeyDWK4dSv7xdNTsp
SRWh7ohsOTweO9t67PTmAd1lM5Zjhxc2ppxaExsgoyU+aEhwCEjsZG8XpmRfbHUb
zGYGR70Jw+SOrPP4L8I1/aNX7qXaZhsqo6KUyx1CdTx+fS7/rHJNABRji7VzXdES
rgjD+OMeElmlo/BzCSQ/PbqU2wqnMd9urLC/D4mUywmDK45cTTqcYLT9OSOkZLSa
e+lUXX2L5H+8WxDvcgTCQNxeVWPHqjAqZeOWbTZL3L18MWD2HPMXdvzxuxKp86Ae
L4ndgo/wMJV3qt4seRk3RRdHfONoY7HqutKucZvcgmIzI8tAvqM2gnvc198GhFcT
ayA8u2HNYE91VP31e+quyDANoCwzAKStWVjBTYtMMcnVfyVNti8zdVxQ9enWf7eY
O0sSa8VZkdCJ5SCPgU0M7nDgroj+GIX/ZqzYOJH6N2J/WgD8IzLP6rq6cl11h0Hy
vPgjYFSsl1MZauvbkl4Rrr2V3YhZldaB5FZKvULCU+JGGt3V+7ZHy+zn2zyMX4eG
Uwr28TprIxpdp3lAEYbx40cr7B50erqCYsF0RQ8c9j31AYtPqtPZJvNFFHkkMbss
xUngDGn7vl/Diqi7Ti2JRC6EWdS0gLW/o8Lg1a6m07VxW1OMydloeLqtd6IcTTp1
Q2+CnNEw0zcJm9YqFfeCQ1b4+pteXVNvQ19F9N2cmwC8lXAaWQVULRqMaqg/lVJ8
iz5mGmitscxONNZGxen/4BEOyh6sf0jeavv7Sh8xqA/HYDKUXDWRGzXrPMDyti2y
o0/nqoTMlQj7TDqRn/R3NGf0yyPSCWC3MC4DkaB5QBqWSSzotGbRuch89wVnwPNh
7Al3j6ZvjVAX69X1qERYMoR38Ouw5Ruez2WMUpFw+xv3COix8xnO7woLJepwmy5X
YH2xVbXuzNGf8HgFLqS5jfHeCVY9FhrxbcpLt1Q0Lq1zQmv15jVYJ7ypu9N5NLji
TLReicg5WG9xk6Le9d2f4p5ZampunVYzqp9/bSD5/mbYCTzfXr5WeHEyYBYRLOqT
WaAShVdQ1UXifscmsGP8XulOBg0QPGa+pE20MKyCgSPUbKxcgUDS+DgxStJSWQPn
UrEC2Ga4OU8tAeBzYEF5hRNP94sC56AS60RLAZSfp3QhRkuI3Wgb0wA7RfB5yXnT
Y8gYajToqswh0RpJDhV80Qzt//+lfiMg0Ke3gCWroo0JXZWW3f0JArnPHsahlYWr
TdPCcjhjzyjXSTNC/EBOZGp7MU6cigirQm2VYQdJLCvt4o898EdNf9nhZSpyU9hZ
SUFDCoWsOVQ6gvaSe/Sak4aAlTOiztEMWZVCEd9yhv3rbVpakvZcxiSJSgD8OKMN
2z7CusVDKPl8bLYQ9/8fKuz/0Gm7y3RS90xfTADbdpGGNp36mPNaWtOQAnSU8jz6
GnZWJe95mmy+9Qzqn7X5W8Rcqdzqscb/+hJUm62GyHn7KUa/yIGxpllzHIBFmrkG
xM7lOBC3mn3S45A2aveXYizhT5qc8CgWOzboI1IG1KjW7BwI8wK3QxcyiKbxSxqj
9fESbxvun3DlPjWfbcCk23BcrwudJZGDpSBm/Jntcly2Pq95HlZ3cISVrYLw2cOO
8IUcFDuuXUT3Voiw9RU+Z1QWUEtkvyOzcCmtFTmQYbaSFzUFVM/PfneT5H5dgXgV
//fzGZgiFGaFZEeeOHkhIdEFhkkPpQ70Uod7DsMe0qYHwef8ZsmbCLgrvM+i1kVm
eDp8XYzZ1qIYjRVzjm4ZvLyDtxiZZB2wHGLz0WmKWqSiNUOzJiVPjrAZvJrN9xm5
Y8NVWsRNJSn3LUiOloEGF4QSwaYCIsp0mJr82l2JjL/+9AYdn5DWBpDRlpRQxZlS
WkZZDa4L8ZyrHavCOhbIQwYAP+xmc61yH/LHuB60mLhyQzPEDvjKxsfiHuFi+EOE
DrGYbILxtD3XxpNmjYC0y2z6HdM7janyAyO9Ds0yW5oHaWtFsijN5jS2JiaMbMSw
0qlH0/+RHYI/fOXN3ty57MQOkJFyIeg13SYWMmnS04BR0WyAzWVSFDtx895ZFG0T
xg+jr8Aj1o6DKSaNYKPE9HfRNq7c28zbtJH5DLociFCyLlXdnM1CX459rcOvl1H8
MAHR+AovcRgQgfu+26kabGhg4FDYFZA+7E8D2mzzvhlTlMJzTFxD9JHQ2VY2DX0R
S619dgBWA+LmTCczLwrP4rl/ZegCPt2h1MFde85+PtOhR+JbjM8zmQPVJmfKPG/S
ZYnqz/Vk1XAZ6uDUCQbxoPTwh2N312kaWGZyUb/gJovNROj7di0x09aJfAGLJm7U
PX0A5vMv+yb8TYdK8PTq9L/9W9oFjxkd55kyFk1NrLqZvXWnQCAGCqVKhIEAoUhy
HduugGWw0sKzsGHAhP3JgF2a1FRLiIi9PXkcGYn4GS56axqNo743ugrwcZBv5k83
907Jro1ZcaFqDT/jJO5Ol9ZV7rD8OFrNq6tF2+aLMP4WrhaG8qxyhNbryyADbYJF
n7F9YP++kmD0rJtOB17BI4mTpTuoEOYHcjLmdggn12kjhgQiWTvYxztXWVbwVl3Q
G01RWikpstD8TfGIvYkvz9xhKrBphd1e4+P5vEkKJZu3MC2hr9idgPEyYg/ZI7P9
aeFs+8jR68dErv9LnB2nEK6dS55KH5BVRN7ysV0gS+wRCNfMTsvfxmuQRy2FMLF6
yzjNdXy8t6saZKOlN2rPtXZon3iwRTQbC2m8x/pARxA9WK/iVZ58pjta6/U/2Ncf
dHh/i8aEvJQEuhbX0iS8QLBilBWWIABCEy6D1eOG0DWt7luaf8/99u5rhrjJNp+N
djFy5iPNoZx1YwDe1muXerSe0xFmh8wiuzKsCX0aIDfsX7xxUdtpQrBJ0Z4hVjvJ
LuoDZyiWS4ey5g3Xi0VoIlzVDvpTGV1fy7FBmrxF9O6IjYXE4WijimsqVhQOz+WH
whBQC13qVTdlrPjE4E51Amgma95iHl4gti7N+mU0EkVxT3T+3H4Aujs8XhVcb63C
qGnpEpV/RyVrdD4NmQ25pD0ASRFh/GqmwUqYWoBhaP1LUQwhcxRBWZ/01VbF9rJD
aRhFXDYrjb0djDDoGMbq/gSWLfoscP1u3pBVLpY8FULTOE6dtXLCd6Pew4gUwUy3
1JNXnvk5og35HByApqwK3nfdmIyViDdyRIoz4ZGAvjMl//eNypqbBJRCH/++Fn4Z
sIDdgNsgBFjFUs37rTgPbzKum/Dv8IjUp91TF0jnEk1hfwPoV15VnhoUNAL9BFeT
jm/8zLua/ELFRl0Ttr4+6tNoWXO/OFcRIVl2rydxTs4eyMHsDiM1K++680HqWLCZ
hM30XYwHN3lvE6zxbuQZhYTwLz2JoVk6soYcni0YxQWZYiXsWe6zNCAzbmc4f1Nz
ifOvYswFq2l8xOk3E+Cygvv9Xm641O4cSSefdwKY9QW7FskVMSx0bxOs56nAmKSg
GpsPWKyPYz2vyNnOyQHXS0wKhM+9QwMPy5W1MaH/pO9H9UNlPINOe3iRX4+oQe/X
SgLRHEhMT9N9HTqDOdfGphzQNsFwdMhOJUYQOYVZNVVHqKIxtP+2+jDWZDHbEPo/
nRJgm+UcoevK6nccbuI5YRGP67Vm9x3+BGjaeVxQq0EUSStf1Ld+xpoW6fQrhKv/
GcJZtD9wLta4sbAvm5doGjQgHRBv8HS9/VpHJoqMo+uN6VUINSSxj4hS/6rtpyQg
4G4vJgH7Uaazve8G1SFC9LYvJe/9GIAXYhDxXsdG7yhE+c/IWPAU71xQSvbXCoF3
ZZYCGhOVhmKYkhyfZZ2CUxWL/UQ2y+NFvSbfW8jvYyjcUPwemsrJ+ORK5l4nT71Q
+FQhlaQc1xJM8ZeBiCB/Q2UFjPGsRAjNfX7BnmYa0qzjZRjbzCjnsoqbxpYkB8VL
cVoPByZt1AHBg649NKNlDIqCQlUnzBQxSWFQkBaFi0oRji8Jm2g0cYLh2Ao0BTkR
kSOv4+TTxoo4rladtds7sSpKp4Qgrcg0jOB3nTHMsMgbggjFaId4JXnwEBBcjwDf
5FRbNXb11pEHwZzNVbYFt77lNYMx+7hFezDEujfQJWqcrvjcKBAyApt21k1tC1pI
ez1wRqlgfQKXKiIYAtbr9j2+JSyu9dKWmISC7n7CwFc01kzRtKDheAvSm/Gogj4R
9czYBe4WcKbzsb6s5yhBReg+30Gkhb6eYT11plIM9CvaKQZ5H4WE8/yvB2Jnq6wj
oYb/zaPkU9BOyYqwvd3o7QEODi3yPGs1pcZMlAKIOE7J5kpHIwN+LjaGmODDmWSa
vyCP0FqgkL9lv0Nbfw7qe67uv9FWQU2Oedwj6e5CXd4Ddmwfgaf/legqtMhzB5RU
X4P9uXqYvSqIZ/rIosmqG/NDcWrSxU3DrrBenLY/IoHcNuyVE+e4arSxYc0CRFDt
oLmshrVar+mji85eIQOlmJIC4l0R1I5zNykj3i7HowbM+aP39KPsWXI7Lcgm9OCb
mpbiQO6VU20SBXdbXsowWac8Zd7HF6ptYycxx6DL2NpsqCH3+nwq1Axm0pyD6872
8FgkdN0edAGcbFDC/aHVG8r6Me/CVZhaBsJxYGEe5OW7Il4T8KOIT+lfKZwuNy3x
450gOTMLN0Buw/FvRXisCeUdX1cANA8jkezHQt271pIUeosU3deIWYILyMnHc/MD
IO2hWgLwaIKhPoHXPgbMIM9oRdkwLe0+0zd8vSgeGG5x6/vXIAKyE7JtppZfGGIa
viGMy1Qg+gtm3RXblSK9j5tX9/HKEn8VAKUfuJUTSQw/82WPNd+jqFldtc3PpgBx
QHxU3TZpMb3KvGMsGusPopUnuWf7OTrv65jGIG38oR5SkYAPsLL2ubK59zpFfGD5
Q4pA8vA3RsnaDckhcnFdi+8EM48E91/J8HY0aeA6nZYkgzwpygfMjQb0QGHK/vdg
OCLhKz+4KHMAzeA75QMyULfBCpujTHCmupqOo7pfcHzQBYsNkNY7lZkJ6JN4bGQA
uGYsc40Dv8FdbfHQ74kQDq/71g5ueUTUrJcqmgkbLBoE2VoqmmvVEXMQ3eUNT//W
mO9176BgaQ7WVz6CXGDQdXCFx9PmaLxfGgavQ6edE0Znm3d3wSbfE2hz3ACpt6Of
i8aSGRNTPENd7OBsd5KUXaKBRTmxmOWy8NNTg+7VL41nII0/Soow858kvQo5NufY
yIKWRk9MgOEs4gTZyMe76ln7MI/WCO0orjpIP9wCgYD/UDLlUkiZGBDztwQ5C4cX
wRADtKyvZNmtJMz6YxVdA+NN2FEEz2Q+akpeNIR9cOh5XiHmrMrPRcf6lI/KlSHi
Cf/Xb9ys8W4xnLWSsArk+fybxjhoarj8/HZoIFlkia7vc+VPzw8s7QosKJGfV9Cy
xhrUQ1+Y0O/zYS4DiPjveo6/8j01zRnwimJaTDL2xPEk7cZAo3krhaV6WOG0x7PI
CMX7Ee2C/V0mmojv8AKMKFWvp0eO2dFciAaVlTMVItbX/wheGizkG+WEMRQOtJYY
sbYMpWrjuw0eGl3NFwqCbpLInWq+3Kf8AwCEZMIofUE8ICXWeKKOTatAgm6BS4a7
KtuCT4t/H6ZL36e7KT52QJ2m3/nMf2/FHIuZfF9fP0rNyPQgkAo0AhwDqFEci6TV
aw2mTopIhEfC/6dEr/3jHpJC+sKyyVL/NvuCREK01VBb+sVIsBoyfiMSZcQTHr/t
R8F2CBGLng4INLqXwy2RmlQ+vx2vXvZaa1LK45SaFXR5fZiGc18vtm3ajeBNSB0H
ez8DVC2AXCRcrnaPc8D11qVzHrwtEEXjHsPMrdIHapMavgQQvSp2pzZ6jTgmej7B
2gYUMvhE2RVVXu9Y+tpnyc5o3FLBaH3t7+yqK8uCquJNP6JrFQrlNsmnSe6wrhV2
7pSVYgRl38PlhLukbtt/YmR4ltvtQk89qwXgkrghJOygDpDJCxkVb8imjwqxznO3
l7sO+UTi5f4AdpvrrsgYPFtwaVR8iCgFUv8V4CBb1fG/Hbvd+fUbt0StohF/Y0B+
FXEbxO4vqe8pWq0SATGFDYUWHtbYLiGSah5xnLlUhfRR1XCodPZ+KtUnFM5EXXup
HEZFf8lIhTXHZriSBa7aDQjynXHA3Hxklhsmf6c3z5PZSz8Qb8AQrFe0/KeNGbcB
4jLjfDOX+tqlKo+QM30ASwG9Aozbd1bX16n6qpATkARTAQSeI8LLT9OXN3EuaY3d
rIX3kxNpUjCy4KOoL1HtBeO9tVzBhwV7aJqfO4T2K8xmBKea2sd8CWSMZPj7i/NK
NzMrjVkd+YSyYabewDjSyxk6effWfq4cosmW3f78Mb13j2c29j/jydIby4XVj0G6
sdL7+u/TF3GqvjfZ9gE+e312akXsXrW+D7ZzCL0cXl8FeEAYTzOtwZMybdE/8vxA
/IkHVpdMm0VZh/Ej/mQU5YSF2f61KRxmbic4Aq1r2hcKdSTEkulbZBDrEBhjj+iV
VgZmdUbDRocYVCloiyBhqKwkptZ3qHqkwYOb74GdttfKHhVMXv8t+U28xVHWKQPh
Uk0qJwyMLsf2R7PA5kadjgIhfSyOuBR0snABdCNDiaNKqKSVBOSo/bTibeZ+Odw2
BjEPCSN0L8c8YB1Vk8b0cIGYC6nus7dyYlrNkzFqqDqLG9SLT4iXPQtihPd3oXQI
szPLMbBpKMfCFKrJy3ShU2jZ+m8ANpy7JTCvskn5BoHW6fPo+89xE+Hb3kRUflKX
19DJDvDwqeUFAXef9fXIZITf2hAQu6J6reqJYSKsCxshjtA5jud15CRygLnH3mKQ
4A46DNK3osKbD5pSCAgSlW9nbs2gYmtFoSKSbMrR5ugu9gvvVBMzO6NxyIrM43jG
79VnOapW5vl9OOOY6lteY94jPekWr1r35ojHuHHgGIfxb8T36DJKVgLmep9VDMul
J+BrslucVF+OrwgWDnEWpUHHAzw983MCFRVfREYZKZCUp5KiZOGbEKT58VxI1Qfh
wpWUA5uEoJE103UjWQqNai5KyBsWHo6dzFbEca82Qsis3usMl+KfWO6yvYFXE0wD
qfOwdfiwrAxLBBe1T5Dn5q+aIayMikIPCjLmQDk3cEL/HuPQQLq/s7kSesNrCDuX
i/SxtPVOK7xH6SU7srAmJKdTMBLoGRwaH2PsLjqHgswAzCMJzsQo8IrhIEa3d5gs
olt55OXqYQFQZPz6hCUnYgk+YPcCvaWg0zTpD3SHgK4N79PlrQOLTccbW7he0FIn
OEeeTrkFpkDRlwu6SQaN+6BpNmDoBPGZDa3wc6x1BI5L7jIuBvZAZOEzmShuxTgy
iWz3/b9KCQ8rJxlqV7TbX9sN99Aj0c9IDEK1Qd7I2IbKPydeeM2yu9Oe24ppY5GO
A6gXAg+L40XyxNY4a+5/WysVn9TzYUxccNfI3mEL9sTw7U8KyFgXiEx+NcJB8BC8
M1DYM7IUCB1IkcWnMa24lfT8YpNLd62Pu3r59KL5qx0c8HjNkOZfi1pNBrE/uI/B
BsYFrW6UDPq1gCZma9jgsLW+koHLUM8Ne10KYhwIqPyAv7hwF9Z1b33n2wcvLQe0
6TGY+GDJq3c5qMlFp4Aq1Uymg5Ywss4PcSxrgXuyNZbwt4oz6cJBQB6nJtoFRnjD
OaisyXse5WiI6u8uGqFyfjbCdf8M1VrNEQkavE0QvpYhnk1aNqzZxmkjbe68lBh/
vZGxELvum58cNTnVrPKb76X3TkY5aIB93hV8jCzHQW7gRT3spBLTf2vnxPsKUSkF
lW0w6k7BRLv4NXdEwlkHxe/t+5AXp6QIovmZPLnwDzhIFrmmAqVueJhnALLyHTR8
elzwOo3B2GucqT7OVI+kMzSR0p5opalDqVNfkXSr0G7g05bGRhLx/FWVQxYbjCYS
sRdTU1jmk1qF86YmXJAqQZrQ4GL13wdh71HtT6qOl8PpCcOhY7/vX0zljt3dd7gV
ZTMtyAbYv47yU3/gj017bhJLb7TtoS4D320flsJiDKcEcQXpPvppcdpWvSw44GNQ
S6ZCZWJTQY7V+MtVFzBtsD0uNndkg7vOrCbdXOLt8mq9jOo6fqLStheWtaiwY9PI
358+OtGvjM19FAioYGvEiWBIefxxv4v+Eu7u5OAD/vrTrk+csVv3PgDW0DT/x53G
n1HHhxoawz3nu6RsWQ0Px18dgJcJmfGlt7qC82kIOF4rHzrC4O5kmITNbiuUp64T
y2oBWmpZJHLTW7Q4JJz0GKLW+QSH7rATjvLA54PzTRDVugWqh2FbFFVuf8BGzSKa
hK8kEenkhl2fb0G+W5HcIXpAKOkKbCn+OtG+5GDx4lb3r3Z7iO5ESUhYohAI9NQo
AZSQj1fHbtjTWTj1ez5QN0bS3X3Tf6fXSxrwAqK85dDkhLynF7VMDQOFCYg4Mpw/
wT1kx83VdB7p7xGaO9c/6Jv5EXFLdX3EFm8eTZN6WpRQdM/vhLozHgmhRFn+ocP0
GeXl4yql/o0jW7AHNnc3Au4kYfnBxzwElLYTYaIr3bu1p2rB4kStOIgWimBRmm7O
goFMGg3nYTAewzUdxgK2iRqbss3zLFV9mzDiXTzAwCcVY4q+v82RXD+lroZbPVae
1aqDAJAWwBtSr6jN6EkN76So2T6agzFXjsvWSsrNVw2+4CwtIVov2RCCTUZob23G
58TEK+s6r1DpiVOakksZ1XX2Rj/0pMhtQIvEOLjzYWUyO6daBWx0qy0erW2x4+br
es+ucrfW9XnEyQAu79lKGUwFbpYXdT25l5ntGvNi3sSf/IxUdJgbglJqbDpE2O7P
4dbwmoNPopAvuvGEiRipHKC3/ANVTaUOXB0i3VeUAflDLgOks3/Nuwk+GRTcjW/v
x6dJC4i2kFvhLGp/ftC/q2Mu+X7gbZpEENUJhKrTW9zGXBUKiGqIiaTxtzdKgzmo
tmciNNp+VcIIaNQGp1VvcsFsUw2gu2TRRtxtZnihviuBH5HPChWIl++9NMMewcn4
76e6kMwzCePyJMqAuxwMss64Eezxbv4FYQPmismuzjldsJtPxIOXmqVhi4RGEkxx
16Gs4eBEwf8wYuKZAKB24ddGzXO00M4QqBl6WfqGFyCpUayNel+PU13nHTWbI5wc
uIF4T0dJ1Xyg7Whki6jR/T4uTwc7hrXsMJ69A1oLxUcOAd2iTIWty2zWJs6dCiVj
6qoZGTfpSvGPKgHxQ5dk8eJ0NwvR1fyrJ2bp6Jo3pHLYju3ezuywFCm+zQGuqbKf
YL7FWXcsPoEtZw2qfSGUngEVxGZlIdARUwhA6/vJM55qJlNRHytVpWJYa+9GJRGB
VS1NunURaRbtLxQG4zOrZDmC+80AWVWYbr4f5O7B4xStIbDY04Hq29J4H6suvhIy
VnPRCXqOY+VUQw4rhL6kr5t/72c0WJvObjwJoRe4dCU/HtaNZylpPXuf53or5dmu
Ajdlp/X7BLFZFb/ggAupn5z3HPXVzoCbySfAgNqya4zecFkWZr0D5tXocT2igukM
wako5PfuvmoWB53vA0Dj4t09yva35AY4T+RoAgyC634BdSjP3hVHqNoCepqpGwDa
ZkSUZDQ3uy/CCgcaSW0OEdie4lpLJZzrwbg+xxCmTSRsHjNCkqEgLcRUnZhRiBlj
3vYepwea9/P0DLFvoxdpUID9QgCNcfcZwWOii41TBqsJlACWR+o3T5UzDtTcbpzv
yrnCV+/v9XaYTw/olGzn4sryidwhvziRMQeKZht6z+JVPfeX5EoEk3Zm5Kaz+Z9R
mBDYoFql1ChsThb6+I4CNvoCzhXCvDD9iK9I/JokgV2FrOkaVrjLImW04m12aYgW
LpCKj26MuxVPKS0CMHs0bhU+9II7Ajg1l1x/9TOL0mUMQgkSlrslvKRNReLpXn3q
aP4A5ff5ehR1TOmDsgYaB+GSQ18M5GVAnLEcmDhGRK2pW6WwLCL95cS77E3mZYe6
8kTotSntODh47/Yxl68Wpbbx0Efj8xdq2dzNwLB55XNXE2zJQ0jWueuDfgKxsJ2r
eqy0NRq6yEN5w/QUMy7HV52r/WHfU1QOlgESI7Fq9wpswsXSpTRITtNr1BPoZHGp
ksx5jlNknJn85ZWUPgQlOQO3yzDy0+Xj0WoyjcUaeOu3JfLviOBSkS5JcyIgx3xH
r/yV/P9beRcw68HZGiq/62+g1hi9rSuIE8dlBiJGox3lmogo0/VM0e4g7dJr6GGz
q3pdyfpWDSEPgjpicE4AW5HzZLq3/ciz1RYKYD1A0P9UT2i9LPBvzgptXAqkFQHW
Gzg265gHunPBk9mYH5TqpA0g4B+ku2bCySuz7vuuaHB3EZi5Y2k1kT5KLBG86Epn
fb4RkGpLvZtDJzwCD0F3dIQ4JJKGqefeM0xYj4+tynrTLoCG8pQXebK9GJSF75k5
eUjyfWBuyJpmh2QHIHJj66M/ZJ/3jhmKi0A/MZqIf8iQcZjvTlhSGrB8xfdYFtJJ
BqoA8OOKythuH5PQS0+NOT2HemIREBmi8tmlcO8nEhxjgAA93WkmZT+HZFeHDgOK
Y2ENwgVrGNjIorumWHkPYQqXBPqxpgdy2scPh7Pi3QpHB/I4LzL675MGoCXcJAA8
gPgSWp5aStZWGqcKeXauZxIIkJT845sKCnyITKu3GgRynW2kPqXhocbqcPJ8nP/c
pdRYdJHXDGEfV4h81WAK/nZGJ8X58vuOn79wXT79LCWqUAymKsRzSAwz6rnaF0wW
PxgeAJhQ8v767pA0W6V7wPeOvcLWoR1ynCw+oAT3Ixs/NX2mJfG4PxUMDyY6utnw
bd9FcYU7GBF46LoFZHs79T1XiWrIWCWPbsHUszWTTeedmbjYUg9f7szy0t7/9hBl
+QOt1wiQaxdwSs1y3bq2wfWEIKWKCN6vDbbep5kj0AaMpwDPD8hP0o08Eq/TM0MT
F6eysmrd5VFUBXbVk/RmxjoqXVOBXqMpxzwoSijGcc0kxa6hFimj5coc8YC+H+0x
qtSwnFb3HrQdNzi88vPWX1Das72wiqVUjGZqx5pX9Q+mUlwEWnrIUPHS7tAH4ViY
PuVpl7X7UGoW5aMyl8IophD8xxojP7p7pemoIkp8givK1UO9vuRa+Sk9QAlvORkS
JEBcr4mi8qILlS6zqTBnG5zT11griLZszTrzWVUE8QO21GsetmRbZxd3CbRW6xrc
x+7B6p/atw8cl1oq4YxKRdgBOcCQskhwolS/QVoD/YXX4OnrOSNDC6OOWxgzUyVj
luf1cigJad5wIDfXjlHv2GQLAX4omoOlc7+ajZb4ZTRnQHsY7caK7bLe3C/WK/mb
L3VwDyfQnRNgdSYN18rJTp0WSHXJ5vBNvjxBL8aSTik8f5tn/E7AjycTP2W185C5
OUeHBbWM4vCAQlOACd00V8eu6zJRCqL/CK2Y3LViSmL9AR6jj8JydFnOeXwcLfxM
YBLtSsX19d37/5ROwDGH2/c5ZBS1cGXkNyuvQlhPYodueXB6sOXnGytDxVeC2XJb
LNi/SQAIyfacbnWKAae/Rt+iHSpoYb5BJ2sEKA9xzCTI5EcZFll8W15ZgqoMsKre
yZbqxvsz/R0VL01zvR4XStjRn2bnt4qQWtZ1btKO9Kn7jENLT31EonVcw4Yr/tLJ
FrPHAd7/t/LSnFUrOiECVFJ19cbT0Os4JKrHvwbbtkcTPkGgb4BtFZ9W7Bjxphpe
1R3YAoNAPUaGGcbqK51hiyFZGwKGursAPOnTSgM3MX3iJ0Z41mSpIoPRw25BToLK
RotRH46H6vSQfrnmc0suM+uJIYZlsgP3nh04btqRWp1t9xnRhtcsQmu74QrVhoNt
AqI9FbS5NskGN5tjEtfm6xTfVghBVi+vJ/4wv9czcbngdTBIhrLFN5lph6dOyxr0
MuLnoR0TW4Y9xJcsWvmrbN1UwS92u5Qeo8RrdmsYQI4wO1EfG7LWWfSRPyUQEeEH
0wpDjIvppVceaFWOXUoV08rubwkRhgTz+6Wcku3Z/SXNXRQa/L37mrQOEjelcTCa
jE1+wjAHEKyW69Ez1bEmruYYv42kpWb0CZWJAYdLNLAy1TrYZXxgXyUfZlIBBdV+
0UV/hsfIw+awTbUxtk1bPvN6RyzlKR0+YEj9BSMMK1k9UphNN+M8PZqXnJuiToJO
mo2Pod4eRPwPVNUZUPY2EWaoEHrmXzwu81x1CUcUbvgTPLO8qv3f3SojFmmW+dyI
V+A2zRBQYHCMmm0cAaFgpApDHuN0ccNGJjVPITF7wY94eZJ+O3h13pQyy4/N4GHi
pThoHHJl+NE3j9/mHu6ncA6sfob3tnv1T2H/d3HqXFCcS5xsoh/eaXkOK/jmvcRp
VbWU/zBRT+SJGmXuzUW0lUuG3EK4r0o/v2xMrStouoch2Iu7R2+HryNDDSMMfMa/
iI647OqNWJ/cmqwNtLAjiYblem3AfLVtyh1OvxUtHcRdhwb8C8zJFwxpBUtlC0cM
D+rovTYs9DQgWOWnB20N0xKd3dYFG8zyiLpfVFOEi+PzMBLJD6LJmIpUZTqLwJUc
9POOEiye2bbgWI6E2alrHNBnZ6WeRbN0T6Z87pCXyTOzTqyGLV6/6tpJ4JAMGoQ5
gR2gLnwp8GqJjB1vh20Zqlb/zy0mCKC8nOGCCrSRQaVt/WfHOnanPfdhcP7odQJX
s2uPK1TVyOEX12xGvuJomXu/t5FK87W4j68wPLjFkK/YQ8tCq7AMeRRXG/lv+WSY
mIWZwbTjH40cJEjkDTs24mAv/asv9WtZ7hA7dB2P6hzOxbqC17/Qrir3Rts/dYOP
VCS9o3iXnkFuCE0U2W39suHp4HwPKpKSuXsnJmmur1ElW2Z96lGALeS60WiPTx3y
fryi5IOOD3+jpjBfrjffhQ02oWgKFhN0318hkUbuI7R11zS3ZNUbmWiY9UscFcUn
E1dfdnt2jSB77B/nK5Gh93Erw0F2xoP/45PIILcuHoXQC95B/KvopxiWNU+AkvRu
7kdY2Ioy1/2myKfZ9NAcrlQkxQn4ECheJaWdjZZOsmn1R4mgtuRjATyFovNn6cqX
Nxbodx+U05mKfLrQN8egs67rmffC7S71ZWkEyhx+6qCFbEoofKWWGU1q5vXIbKLh
3uQ962qQPnp9qSDKHTh7yUv8iqzCj+7Q2NnpNgd0ExcbxGtJcCaZfyfIu5E4gQkZ
XPxKM0TcwLSextTSJIz6YHtu/6qTjMmcPX3PiaEnAE5dFBkt79Aw2TJO4r+eESiw
bPfg67/kUleqrChsRGuClqI629PTEJj/AtQgognCEJSxHP4Ua4Z7ReFveaTXVswi
zdfZeqaR5agu8RXMu8v9kXvew95CpZHsrWF25bGUphIymOsLvpMaaC7a2/DRmIWW
3HL4IP2Td0yh3ZK+D5Bf0s3Z119rGRWK8cxJiwVa0ie5dEyyA20Q4yytRrhH+wPK
3HqkO1dhztIJXM1aKwAz3I9xJj6NsNwzcOYxPtveQdr/slPZP7AbjRYNOECjXY59
4FBK9R3wajDP3p1hCP4IVTQ6gSzLmLdAXG3jpYjvNvaEnef5aRJJ85M84aOEx3rZ
/yByd4qAUyf1iq2vVTJmmd9S1xW9DZxI99J2gTZgy4/rqBWBq+PSpu3dsPT3HApE
A3XjAfW+mmAL8eA9DrOWalVWFkrgSKe8wJhqEMtRB2UZo83ziBnylsbZnSiutmG1
SOLXRo9ObAxf4H2fJ3OYU+W0WB/yD+dZMRGev0KyJA6f9wf2NeklQB39iYZndO/k
o1C2A+qt0SjMdbPRUQ3KHmNQGIp9mxOTztnPU3D5HQsxbEk4kuf4I9EJcog1A4qu
vmjqh8XijGg7CMlLtq7kIAOUsqBOyk7byoU6u5zcMZoQ43PLnc4NSyrgVdtdKEeV
+NQNrr+Jznnj3EJuEpFo3r+Vzkb8/Rrfc64CCZ9CfbLe9GcEhbLuJVv44MR4yvre
2KoPf0lffwXaUJ2qB3kiHQJhJP3hrrCoJ8r9E5K1KKBuRALwqXAORGpFikKmjW/A
sXCD3xoHmhGk3KCWYdDFM1B148H28+TTN/G1adO5GSFjwBHSshrdf6F/sUR6eAOQ
D1ALyNcEndd4Uwif3quUoskRvY/Wp5/MObJ9icrqrr8xFhVODaJpj/SO4Mny0UwT
Z9Hzk8LsFuEePOI50fEvHqIwtpTSQhR5E/xzGwA8kH+8S/owlfoSgv5lDSIjVRAs
gFNaNkhxGM5zt87pHMW6zIjgLSDpfjxwEbaaJJ2k2mSq8KIWVA0z6cL1Fhn6BaJ0
nrjgU27DNoJdKCf8Q7Gh1URO/Je9xhnbbcxUXD2wkIPkBfnzl5krbvqDt28deOLs
htlYguKWl67Jm/4+LzBvYmwsAhmXD/QFnmBI3FA9ZDqGJwmv/GlotrG5kh6Szexn
wXCkGH83ZRNbyrLxDOJXF+6AzdVZNZ5rBklKFCegjh8VxRKd1/WSIC3PuhOKRehJ
NcPloBTRiHDvOz9nteposL4Ywz9pyT6fSktW1g2KBr5ZjyDcNQbdHZmabEm7+ULL
rjWlQ9yX80l7TvxOGG8wo/Emk/KlevgLoIHHJ7Bg21I7WEnde9nmNhCA+oSonSOc
XAm/mHbGXQ6z8tSWMA4nxc8BcgzkBrCnEs2bi9u4FDJki3jDrOFpjr8qO9iqutLr
27kx7BuX1rWt1NN7gFJSaFPMpq9HdiZCBQxheOFlCbyfZs2sOrUi8M1w7pbgn6nB
DJ187XuKTgcO71Xt/2CPDDxv98EO2d/KWxDg79SqWY77RxIJKGvhWabJGVM8JU00
8BXS2nklZBoDdYma23TlgrDIOD+KbUE+DsLtjDo8hru8J9o+pBvon5NhIWyIEay5
5eaeXzdy0HN7E2BZYFvVT0nZz8t9hksySMpTfcMrfOJrctKWmVdUmrJ9K6KokrF0
pZqjtzJlEK4cjlShcnW2hMSmU+iSbD3/jqLr2xqmr1AEJXDs0XVoTqT9xjq5Wun2
64SI35pLwRzLAXoj0bDbjU6A4eltwivssF6ntZlZTtQiiC/JLrLtycW5hMOeX/tK
cS9ZbDgj8/cAKzr9NCqEdRZorpucIr5LmNLaaZH1ft8nXiV8CtCK2YdVLnA1j2TG
cO8sebtcooFcrcIsxpyVpm3NGnIhWIKW19h64LH283ZKoAlRmzUmtLGdSWPREir6
PcMzX8Os2nP9ZffW6e4odHEy8td6uFCHIjaIG/WF2B7jm1hCtnxl9BBcAftVRrXw
BiRzTx36MiOUnELpWvaoSvmTDYkqm2I+uu6tymDzFWfwuXuhoL3kJgLUKFzNxw4B
t6ORruaVVTOsdBryq9RIl84QAf0DnkihEmAjmJA63ObMw5z7fBxJ3AB7C0KaCBft
aOdpH2vdjovxVJAbRGEcT07a0C9osE8EbL8pc2KvvdsNKxXWPdVeG0JIe/tbabTJ
9QkAXyYFYMd6YuRbEWpVip2yO5MmuQigpv7YF8RU/4Q1mCklo8E1Gd7VFWgRMsgW
c44p0H96IjKpWGNb6dmUtN07RwijedEjEhR+45MGnT+NsvWZ2ioImMRQJSAgiJXV
52sIfgoejU/KmHayUcbuTZiJ0APU2dretSVpD43Va9bZkDnxiEt0fYIGulJCvhI1
SjAoLkBIvcpwk13/ZUTPp20MzMNcv170x3SQXgsRMeRCGV0sNT1qqfSZ66f7xNbR
w1UsscOl4INu0cxS+mRHTTDTl+P4UKuoGb0VZ+zCIfHFn30m5NfQFGBwuGRbtpou
/anbL7bZMi9J7Jty8A11AtxYs/8MzrIunt5U76xV24Y7REjgKOJN9gaRTXSA3h7+
ghvhXNrt/wu5YDUdLPbknhuwro4VPBCmKtVVhrHsH6jfs4yroknyUBt/4DcJoBk/
jDCv0bu3ThEYsFYkR5w5qDETN2aNN/Dt0xtEVWn9Y+yvB4HBqgJVLInne5ybbuDC
jeNiTRnxYoNItRWO5fPMNLaicUo17wDCp2vMVOnPVkbta3uR9xw6pXtcY1Ls5aML
wCLDORW3/E0/8fhiBZcwYxX2Re8sEyejrNQUZemgKp2aU8lvFpnm3DBHiEUvquUB
Q75CS7Pll7AOHVs4NRiw6bWW4/TXcFAeiIskIeKi5Bvkx853Ooc2xJftc0XZerjS
0n0F8C9pR4b5yzBrzL2qnt87TIY3WcNhif5uZc//EXg1QeDx1juRmsRiJtqHShF9
xZbNv/7ipgWN9KFTHs57xsfKxChJaJyOl8R8Akm6Uhm/+MlA+23hJ376o/wDXSwx
jHUTdXbQbZXsq89KM7X3gzb+N1Y0t5Uk//Xvg4eDFYWmpbm9+Nox4ys57pZ9mMLl
sEqiEJoDpXRLKgXkrDGDeenq2N5eLSD2TmX7wWa5rZwnkjTXZX38QfeyJRLi1CcW
6f6KKKHgHeA3X2uO+BpbN2mXz7zkboav0OeJnV2KUhWn8P9OcB763t5T7xlCE0/f
t1YNyTwg7WqrdjVRIPEGcQgTtQpfB7+X+xMWRJ6wnNpWpKz5jVF0OYMjj4dlDKI3
55LH+cCTqBFJQzLyO4sAXTUutTDz6anEuXwV4R/84qLRXSKR2KiqscuXFecr4H2W
XEPa8ky7VYN1FxudevAZQdP9sOh/1KW2BvBL5o5/ePVzxqvjX/QG7H2dBjIjv9+b
2F3WNqnSEmD8oUIVXAi6PHshYjBAYS3Zn7EDfyVTBLfF38mfe5RFjz60xii5EHjD
uWZEzVIeKA2wZ2QqbtuzJu3bIPzme20lwTpFu6lfEBwvnuvd2qlHvWgCM5hCWpdD
ZAUHVVVTmBgqwr4pHYrpufBTPCzDyl6Mlij3mncLCXvV6bVxT1L38Dwpx1KdVXol
aRN42HqDq5SXMLIwXdiogEuF6upJv2JX8gva/WQD3CuSdFY0fQfLm4KsITr6Z40r
N1l+4/WpgzVf3M0YPEjdLdShoEBPXrlGmm6GQDuxB27RjBxbH13oNJ2xaI8DdVmJ
TNXWxabsZV6OxuJKdEAe4l9ie05upnxaEWAhP0/ma6i+bP7+1EV7oakXMPcW9p4k
0xxunE8P+mjQ4Jbk7Y1cQMiVWD8/L7G23rq0iJHz8oThrL+6SCA3v9Cv8P9sRklG
ELQ5nLAtwgp+H7RlIwhD2DkCVFjUF0R003QyT8rjgnbyVth4w+qJjw/iTyzR5mvO
ytCxqOgR5hrjS+hIqSOiv31jYyKEP+LxiyoxjXbNFIhgytI6PZS1ncpDAHyhcokN
/r65RBGIBpQqokssSl7E1/OppoeDWN8MoecjazZVoVtqI/lajLEWL4wTdWosQZ/m
6Rvp4ZYeSel0ZlALgljC00LPZxdU2UU8kV0lbrmLYHUgm1GoNED+55R7hk1tAvEB
o2AhkwlLUS21YLw4Ta93PJdhBVGTHynbfu+VTooX0uB669Dj7TsP92vqOscqhXTs
TS01EeZnSBwYjysOwoCzX+L86/a0BtTVTlSHUErXcFlOxXyWEjONLdmmJodxTgWv
Nn2fTvGRjdS976jdZScDoGqZuKVq/pNktg+4e0ET5+uZr8JuY2vcoMBz2yIFfbhe
0YMsFtvdYjsaapHpLutGOrxeOjkCqj9zvwTWyrPn8Vhe0+MXBHbTDyGt0tsZCEoe
TGztMQhOpQVF06hIXkIPQyOpU/uaL2WP1CCB6ixteHN3bgx3ZsJ+ZjLasOvjup1M
ihlWXNQ9s5Qg4lyYbhC5fH0Q29pBaVUmLpwGVofw3ZgKiiQ+1QKIod/9QuPnXAlJ
0tbGmpOPh69Dcxk+0YECFQSYygmkQPY+J8ZQwASV4W6oKGYfI1whEgci503rJMOP
2y921kTGJglzygbuotMdscnfnvMD3rY0BAIKqNsTv0r8V9pUHNtvwerrRUO46GtW
PyG0UqoYcYLxfLZ/T4Wx9H0eVv7xcz7LSnSOkiOarNh+dpc6xVtFjHFuL2mlq61r
10kvxFIvKU7Xe3tAAo6XOdJyoJO7JP/wqpNRfOXAU2mSHJ626OnNIV2PrrDDwPFm
KDeYUjKiakAVKGRwxgoVj8MzLVdjIgfweRaUHUqlRKJx+3I6kv/EMx4H6+YK2bk/
I8purhaFBiUq8SjbPTiX8Y+Ry6oaBYyyNgMNrWHSQr3NshoTGv2jwYD5X7V4hZ5c
Zjbzxo4/GUKQnG4go3/4ZuiEbPIoaBjrhd1UKnK6UL6bXfOnImScgLiU+w1rJDnW
5vMXGk+gQ/GrhsgPmdnZA7jaVnd4gisRObO3enpNXJbUV8z1OR8+/itxHVBBhX5l
NtA/A2cgH1ksxQiqR+MxYbGovWLaXbjAqKUoPsLmvx8bYdDkdDSpl6ufsCTc04gw
y8STbpFRnF2P3Y9QO7VZlSSCH3k/EeKTgXh/JxBu/IVQqd5OkKJLkuEzXlXtuvB3
57DRrReOBT9NgYHhMNvpTegdQ0PnF6C9zZYjtqFhy3Yvk9jUlvRt3BuYa4XTku+Y
v9w2wI7REByPvpGz9ZcE/ojqMIolkAHMFAx+TS7hTqPGGgml9kaIUPZ0/kGVX96T
ZVA5lWhbMO75Y9XfHZY1ShkfEalVRNNc8pRz8fBS1irrdK7zR8iNNGdBdUdrhTbW
E43W+31XNhkwniwkK08DKyOgSGhGhEouJPKWUfkR8GJ3aEFXAALuKwPkWW3P2kAJ
yKOP5GTYBz62cDsV4Ml7x3fgDjv4opQiHLxIHemEL0ukA/WO8nWabX+q7RVCdnLi
H3t8/a+XMPlQJMWqhUpLvYSY17pBirjzdXLDsYHHXl0axKbXkE7ThHzdAbvBBMgV
eLoJx9sPeUixgdOc+8OZLaj9KtnnuXv6Cle3rdpVFLhUovdV86IhEmrzxGyIXw2E
+FQXDd8zIpq2zvbkvueWYj4kLpXKvZMEL+gK2mWN7KMV4nCoSwHSdlYOVXfGXpdt
9QhuPBW8YtRnvUPqwD8LijH0dsZERNdPwsJcUyw4HA7AYIyqZm1pUy63PjHC+L5s
pc6HeeiP7iGKKIkZIagOquYyxXT2Xpoxqn1kPLww/7FDqUAD4uobmkEKm+AY18oW
zhPtuuKsGs5rIVuCpjlOh2UdeVDsdxQbAlDj5xSFzOUYVa6k6BW0bC4L+z2bm6TS
XSNB4E+nNGQbAxNjABakt5xSTnYbojWvUVYMPqD1tniNlsJZtMWYejnzDlfvlDIL
d8At+t8dltddhxku89o+rXYLBweEU+o0rIBflocNXWjw2emfGyInFfCpIu4HVXhW
7yv0WGeDzwGc5TeFXVXLa9RwiCof5EsJdb0uwKTJ42D5sS6CgLdNMcTyJYpVNb+Z
QrtyFKYHi93N2rjGVClRlGCoapSNrm08UKVXzrmhME/uwIZNCdzMGgO9Sa9gaKeR
pFxV8X7V8ikDhnut2AWtCiWzqrI6kbo76xIfnQNOClnBsLui7k9/KjsQvwd6Go0w
WVq2y89RHrHC6DboQm42CobYEuUc7SVmjLralSfnIEd50YFaMqQ8KUwl+I76FoiA
U9mkUhac6BZ9JzfaxnHaaCTlcFifqvGW6SFyNBG6BNdJ1R/zvjT3pffTl8k/JU2Z
FSqGSxmG8GWLdpUWrJbHbFTubzhJHHMeibihzn5aTXpmaC6sT+iCbSwWtyDdaDeI
MQ+EfMZSgHXrOBwO+rg5xBigoowTD1wCN9so+d8F6TfK08v9G7Ivx810ffUDPx2X
+bsZ0VbaJb9RhVV0R7Q/uEMTl0LTVq5HwEMEIzKbEERsBn9EmqPU6HEQLbp40ssA
7vEwLqbO1anrDoQIX2Vd4URCDt5ZJc3CJ1tg7eNvNMOVM0lbgyxme0ZQaCu+vxQL
DiNRzTbw9hZfwNOE7x/PE1pwlJOYj1gR2X4u3qV1VnLRB6Gzm1Q6cpUks0fpn69v
ozJ7gFYbUlte0kaYGjP0a0cma3Pxfk33gHxtdy9z6jPZv3r63LedH7gDb9igG1eT
9VC4DDgo/iqu7ryhuaDZtt//6ActVR+Sm96vbtMT/8ceT/mc7ONZ1w03Mn+4UjSy
qtKHD+Weu/p9scRinCGbDJVv9ojzH/X6DmAVnEUn64tWSXaeDaOloqY4zvIIOPcS
/q10joIHh78ZzmopmKuiv/dGMjm3bV+lRJyu281k4RAxjLYzxP67VA08Ll3jKCqA
TM4gzSK6zmHVJE9wrNtKJX2UkNkGTFQMCpotsDW30h/5Itqbn4Q0yQWBAc8penMd
u67Ji7hRRDlMqUxwXwPUtw19LPbXUuv7452gSauDNQQKUbar8JkgqDOkskxPEG8w
s2KIkBE7aka32jbFs5Pe9APKPbHT9uqpjZJBNdIjEoZYlo4o+mutAKu8IByGV4cM
DRGDTdTF2fMyybbFG2AUJzANso1acg4VZDKxVSf4SCRvEZvmdEdPbOTP4FidDXaW
7UmOAvY5DbY1o7loWbU+dJV5Zk58k6nOjZi19Ts4X9uFV3yavQrC27KFD26RrP3u
4o6uVI71GHgf3EDlwkRq7PVx4MRV8pWKzXqSPyd2086BTp4KELxD4yuGOHO6vnHQ
5RYDjHcnqYJsDfx75APyqD3NFX71fB3CVRy9r5wZzHwX5DoeU9K6Xw0eiBVIrgMq
RUR14q1/OoAgXDM1yu5FnbcfSu22xTjOyQMZGL9qOacqHBEhDY7J3euvvHxAIrtu
MopB+JY8+Eo7007w62xfgUkSVkm/ORQXc844O4ERIhqDfP9XfxGamddbrerBND/q
DFdvwGItPjg2XsWTpdPPfuObY2Z0ET1jToep0p7zLaLQBHSMacu6eXUUCtoR5DhS
+SMr86fYRsQkanLwFYxCvaD1rNl+6A6n4EdYoQ7U4l2IPK6dacejp1Re6sT14CHk
eXcWR/TdHMZEfUBOxZjIoX23PirNMjPZ6NFj9YEERCM1Hbajv2rYE02MyAkhfyrd
qnzZ60D+5sWuoFaofIUoCRJg33swvvRgcaATrPrxtJJyHpNspPrSdPcGmX6JNRQJ
hcxDeZTyF9xPK/v55HoJIjgUD0MA1d6EX1zqFpz5mhuAFX/Wj6AuIra+6alVsGyU
pEp3b09Ui86yuVnl6yY7u25koZjzWsfmWRxrKQI65PE6OZXjP8Oq4LVy/xZglXVP
XoQ0LUwWIb0h92Z2Z5RVlwvs1EzYu3nuT7BzqXETaCzhDMuaVYbr0iismDyjwDpK
V8vqcvZYEpK/MhWKGyzzNWrNHLHk0eCue0/r/j5DxgVD+9JYmB9J0EjFB9teixTN
b66ELnYnBJFjTE6OP0xza2Zmeqv0unhGnmrrjJaoq6eseWEXPuTSYjVSeqv01O6j
4xgj6kFpSvSNMpvhRQAt9gMhAmMRQg7TAIeTjOYQU/+/oAj8fitsZLVXVNmWBC4A
wE+dcU90ZFEkpbXGK9iQ+U70apenIq1AwWWVkv8+xSdvVeEXmVPw3vxmuFQhVDDJ
1h/dDpv8aGP3eLUa/FIQ85n3GJoU16IRi8fSbBVal+RcfpLvArIhmfnk67xamc0X
iQiIIvwQG6uUPf25TFa7ln2Yp2cLEXXYgkADjBXBwb6qhOc7Nz8XsMAkpIOyjha+
ffMXjO0oJRDpV9Xsb1WY87XbfI39pzisX57aPhE1t6AhSyvWNDEXCkpvvDPuNk7s
keKq5iK8XmIa0uHWd6yGs6nRTg5t254uDqPPQ21wr5VF4ntChyoC7o+DVAK7Cl8A
8Rt7rrU2V8tbLP5Lrza/2ucazqakOvC7kNaHnoHI48zfloNTPJSlV+DXt/neNrEr
nYhUu5/5e+OkEO5NtErp65Lykne7I57ta2f1k+15KeMoLa1CkUMkAIgyN5VZatto
mGnfyJmWU9+U1FI+Xp6cxEE9bq7C6chj+riLz3G7Qny6KnZxBqR1labrHJ6HRwql
HO0gfzY4LmtPqydNcs+JJ7JBX+BUG/L0zOc7O1kAm7TZoWcPUx1ZJhkkWh9xLQYy
4wPQN/VtLCiJtGL/nZMCqKVwTjPuspO5lFqjrWwo1R6lH1ruukUZmxmxpz9+aFPh
iZ7A+wUYn8HUCIzAs0ElRtyC51QVkhk9DVJbi1xiAJSkG/98AAv1aWFLlDQQT1mH
S73dbv+1pruCkaw7Aa2YalDj79v5aiCOtmjjDMclUNGGB+CjCIJGokG7Q7rgRoZU
l63sp2hnazQYmUxltJcExD/Z9anJGVxLOde380XhT/5zLpusgE7lJEmc63r005SG
JnB/yszkzQ542PPyPVeOvgmd/azESjkNWZ6jInaUlcvSi5RtlL+5MPpMiCozEBZi
B13QsQVZc04eiQ+MuuFt1RCt20NV8d0LCYMMVKilfvjs4hhkHnBQOTkha4tc4kvc
mu4+JacS3CMvWmvWjjxMnwBW1XqfRhFD4BYF9T2X3zg6CeSGkyaGXsto+o7li0Q2
mMyeT9b1CBG0sZGTB1HQ1B3JG0ZP+D4Fy/RWGJ+PLXk7Zo4nQpmrbVeGdsbqsv11
A4LCfBK7PIuIS1f8qEGUqSxId22jTcCplisCgw4nhbvyUhIjazp14PmRPkbZlVna
+59V4JrBImxuiIuE1r/iZqEeW1owsmm3BbOZ1oaEnsmUiywPcDVxgRNzTMImECdT
upjteP+LnGlrDrD+6rJWTRWZTkCjvfbplGbeWVArN0mb31HI+jh2MYoFucGRZGxM
Fw6ntKkvby+Z67dJLs6uU5LScXIPQqwn++oxAgatjNZwoNT8QKNymK8qV5AQBxNo
t7uEMSbRgX+ovOlNrARtxoY5IsZc0ZyqUyHHgGty0L4LwdfSFcns1XS4wB02Ko2c
3dKvCC3Z6syy5EnolP7KoUZiY967GMG0IiRBRdG5yHCGI+fnaIc0V4ygLm5yMjAU
LJDdxJUciPPcXeuUpUyu+JCpWqLFjJN7Lp2FRZqZLttKQlLLfWnv7CfcaLkGU4Vy
UkSXqZDIBSMF+I+W9Tu3EB0gE9SHC16jsRE3VmcGCD4M5rm7khBDRtrq2g7X5fE5
R+eL5QY/adpb+rlSCUbjduLq6H0xyHuXDkfWtV5RsqBomG7szD35qiIXMP/dB0gE
XazIUhRAUoGLjO0ODrFfsqPRyxJFuhzw4sg5vnJLV/cwizRzlajOzJJeaHoTo7IL
c4InEkkCflteMtjgNMiFK1+LEiP07xuRWSS0D4kYZ36j3lrzBXKOxC7vZEs52ujP
/Y8jTSeqf0LtbsLwkQKBBLF1/61v+VoXISHkqzDLlhS4r/oLBvuyG9dLsfg4J3ku
ILZqllJ/TpYoYEi4VR0VlKo2rXLsne04bjgcnHFyljNigqMrRvD61edmKbxKyslH
zQtN8XBMySx4WFv5LO4bWMmyTsomEmkPaeNKo5yO4FwIxYvy+DNUF3FqXVCNbhbK
JzR+Fdp/slm0BwXmTKlUGH+NnAiAUWuAE8/AORaqG7nYJiZyO4CYeVSnBfHk3Ks3
S4U1MXYx8Y1P7QAamPw7p+SVyFPOsyk2/Mae485UR5lZSr5xV7BzY9WZ57Wc3di8
hnNZ8U9sMxEBKJmNmw3SIpBnCv8a4MmaCPhRAHKoYoUiU7X+WZlzGn/cKiy+zQih
IMR0K7+fxakPYh5NVdSNcgp12iZF+BDgL8vtiWwQlggDBZw3nbI4SOsMrkOmRRim
Oty3LZMNtuJ+D1rJjDojD8DtEu82sziPQ5xm5UchBgCnU4KR+UdEXin30GMjhZdf
HTPqXK7WbTQM9jpMJJDMqYEBI2OngU7ujEggo403TTlVmy3YE/eVs+n1miJPeI/4
LuS6ak3x3KHccRDdITu5tLJI9XaXqSSKfOQujoBGDKTTwB9bl9nEjiSldsg7T982
MViDrsgKrNYKxZ1Tnk5PjWvkfKz9eu4n04TP2PPT9833DbMGnv3cpwRZbVLs7s0o
arvQyn72KjBCaf8bjzRLeYRJ6AE9WwF1TC7qaP6ZwnN2TqhKcRb6FHIHqzd/TJ38
jnKSc8807NKgVtNix3RkAvhlLRLCV8tEuoOzeOvCyXxkCvwrxWXM6P2+l7b5PxyL
g4+Lxs1W2dqt0ETbyhX/Xg0GHFsFoImhLz9J3Goi5oqK58L+z1oSrqRJ16STBj/G
yDp+gjnH7jTBF6jW9KURutRcQB1X1ldrYToOFJuj+PtpX4vJ710dY0R8c15qEwBd
EjIsf8JdSdZBhwEMLSfK5e+7pwURK6RLO3okuJ69KFLVniS+IQA8BBhxDnNyUb4b
ydJTfqF8lL4BRFToNEyfON87V3EPOYhyjsLzph7WAVEKSxwqosEBVyPeZUzZFurl
+4nUAmXqrnoDxyIuE8ewRFtJkO2P+TOBbJwTx1wmXs8H10VvqFHJaqlmhfLjz2me
RNZXd1ec46n49FhOchr5abCLFfQCRsipvWiaVJhr9ZAqtGePAMYRlvTw6cuoka7z
cegvBOXnkVKr6Scc99TRdp4hI+TXoPBhxyNnMOa7qcvnaYJgnuvQ75ol/4nU61k1
nMzf7f4O4EwJDatRnJ2mpryHgI9srnkpx4YL3JXcsaDDqibH4SumBfWPtXPNHiSv
1TyIE3qIh0ViGTo7aBofOjpYz8CPa4hsVzhvxbEI9IN8wJ/LJDVUA08/S/u3qvtH
dsOI8MRlHWx+rTxt4gp88zG6TAwf6xSVZnojEs5XDNzQxKRpWlOzZxHRCnOyKPsQ
lKNWbrIkxPbcm8MEeuetE7OZqvt2gZcRVChfAAnoQZHTwdvLy9xyeKQAsxSt2+t9
5dQRrRohavExtbz2Pl4nzW5nuGkfXkWjPKGN7Afo37ts5ArqMUwFbDmHuB7N6S+q
FMKCaYUu4oBI35IeKkWmAw83785176FhbUWf+O4YjBljKYgNSZu+kjpxEP8XNnyM
/KkZ2XDbAVi3YP2ho8bYPWnAIW58XEE9p2nr5WDEq7aZgboKnInixKAi4EGwZWNc
OiYkNyE32QyvKevRITEGoWVtG0pbes/u64TJ4kZZntvheL75FI0g5pGxH0z2VNhR
IIKLOzowiEgTShaBcChjnfzsJsK92IIKzTXZtdBqz8VlNkQqoN1idlrD6ZKj1vf4
O5MBT27wpE8ms2Kb3ir+6E0fkTcL+l8JmghVCYn8M6rmHgt9Vb7WCkn1yEMn3DB9
9UgVVvHgo92RZUBA5sij886Bu/T9LK1v9IsWcoRcMsLdOc0Bjcbgg3uO84e+onrz
ntxd8JnYDGPk9b/sf/ffj5WN5VKCVRNEigTR32Y8o4Q2fMwpXv1GAXEBP+P64DWs
016rj2h2tfOMgNuz15IBjGXloOlUSq6l0021+91QjbRjKF0tKXM7XsV70Q9soN7r
miPUMYQUTILsYIXN5+j48hLMbUMbI7Ikm2vzXMNm59CppDzyb/DD+m8h4VH6Xzdq
x8BBPjHMvqR3o4zjfyusnXMVLPPY/CCIlonAi/mSQIWBwIn9CEGiohx9ZlKEy/AS
PtNkqo2Y44fXvjpIg/VyhsA6GpdLyAnflA9W+RyBUp3UpbeyjJNTfw6vWuCANnBa
VnFpLPWn77HONLaB7QTy/eOURXLudLM4sweqHi8BSTXRVVHJceveYB6xwQ2IHunv
fmlJdyiOlJADMIHvgqjaJ6/K5pLD5NrE3m2dfrjN1k6GPSqElEJrLZrGKqY38erl
r6ssj/7o977GwyDfrfITXTBY5agL4MZtbBYT9rfNdS8ymkX1xuQfNz9oPZ1cJRXW
DtcnuHvNeoDH/kHM/aHk+mWZJoolkihIcjDYY5XVRNrbqisxsjH1aEvY3UtKPne7
9EADvHVmJjWZDF4ytJIUFglEPu+THWz6VTsPE1JEG2+mvU4NYdZkGtGH2kDazVT4
a0ko1gvL09zxPOmJ7cDlW6gRbgVyPrMyTqmAYoqv4kA5UiRFU58tu90ln2uRFbjK
u/pc9WDSwKNjer/hZasznkrZ9TAumtp0STeNMACyZZ5mfXWPcy1ejQr1t47x8RLl
ZoRFN7n5Hyr+cD5oC4OWjy9Rfztdbx3t4VLmQVaBxcxqEJBhRx/xYa8ZFcA7qJbp
SXYwGXzzdoeTE0QXRUZxE9tN3crbXH7GcoqCv5egpbcUkj92iWHyCD5ZRvTnmaph
vX9qTowsFPbJqWSmKGyus7YQUxmoFnmLkJdAm3CCTHjhes4VXdVo6yUKlK5ENISB
7fhFhKDdL2fHvv+TJM4dujafzJZL+0NKIKqBo3akVJphYx/swO094I76bfCrpz26
IvgWwbcNjgKa47IJbymkp2a6baZOSBGuJkFhm0k9QieJcdOU0+VRHi9lN3HaocRh
AHScnHe6osXges+GaUlgLYZplFXmuzgdbYrONvtVJP2IeXyF/5BQKYiFMOThOLZ5
W9aSea6Al4zCOz9rQuZnowSnKZrczl+0xPe0qu+KKsWS/hQCxC33zxPYW2s129YX
ycEWPDUlQn54Mga8yMVhOnwjJEbEwqVvYbFfHkdljzK7ZjQQ/qpeLsqpnVk3L+rK
Kp05tqxDZL5Hd9DDSKyFhQ8l0/byMWj1HvNs7AD/H765XV2DE80h5+ar2gsp6D1h
bOWAiiSDA5TC4XP/pTnLKWcPOyaLsieEQ7SRQ0PQMbk0dYCrEZvxS1hHHp0tHLi2
3q0n1OIhMEFS/X2QoW8DIoY7QfdSrCsnC9dByeBsb2JyYfb19nv/YgpsFFL9LCPf
IFrB93vSQcHBnR9PiqLRAFCJcrzibuFafYXS42tfrCNqWQcWhSRu8JQwcc8r8etl
P2mKxRmqAPppQUTixPnY+Irf+FqezJ+MJq6XiWc+Wy7hjh7LB1a/MmMygcZ2CW/W
S9NmEDNther4nfB3nr98BZGFfW4jJdUINk55IpD37v8=
`pragma protect end_protected
